magic
tech scmos
timestamp 1732104633
<< nwell >>
rect -818 277 -695 300
rect -689 277 -590 300
rect -818 254 -794 277
rect -719 265 -695 277
rect -614 254 -590 277
rect -582 265 -483 288
rect -507 242 -483 265
rect -431 265 -332 288
rect -431 242 -407 265
rect -322 254 -298 289
rect -269 265 -170 288
rect -163 265 -64 288
rect -194 242 -170 265
rect -88 242 -64 265
rect -751 194 -716 218
rect -682 194 -644 218
rect -744 164 -708 188
rect -672 164 -636 188
rect -574 182 -539 206
rect -505 182 -467 206
rect -390 182 -355 206
rect -321 182 -283 206
rect -208 182 -173 206
rect -139 182 -101 206
rect -68 192 31 215
rect -743 123 -719 158
rect -671 123 -647 158
rect -567 152 -531 176
rect -495 152 -459 176
rect -383 152 -347 176
rect -311 152 -275 176
rect -201 152 -165 176
rect -129 152 -93 176
rect 7 169 31 192
rect -676 83 -652 117
rect -646 83 -622 117
rect -566 111 -542 146
rect -494 111 -470 146
rect -382 111 -358 146
rect -310 111 -286 146
rect -200 111 -176 146
rect -128 111 -104 146
rect -78 114 21 137
rect -499 71 -475 105
rect -469 71 -445 105
rect -315 71 -291 105
rect -285 71 -261 105
rect -133 71 -109 105
rect -103 71 -79 105
rect -3 91 21 114
rect -800 4 -688 38
rect -652 1 -565 35
rect -471 1 -436 25
rect -430 9 -364 43
rect -54 36 45 59
rect 55 36 79 71
rect -287 1 -252 25
rect -867 -44 -843 -9
rect -833 -44 -746 -10
rect -705 -36 -661 -2
rect -487 -40 -443 -6
rect -303 -40 -259 -6
rect -208 -13 -174 31
rect -105 1 -70 25
rect -54 13 -30 36
rect -121 -40 -77 -6
rect -817 -144 -783 -100
rect -742 -121 -655 -87
rect -649 -110 -583 -76
rect -564 -85 -498 -51
rect -380 -82 -314 -48
rect -65 -51 34 -28
rect 10 -74 34 -51
rect -473 -121 -386 -87
rect -227 -104 -128 -81
rect -227 -127 -203 -104
rect 10 -141 34 -118
rect -846 -179 -747 -156
rect -846 -202 -822 -179
rect -766 -232 -731 -208
rect -602 -210 -568 -164
rect -129 -178 -94 -154
rect -65 -164 34 -141
<< ntransistor >>
rect -781 264 -779 269
rect -757 264 -755 269
rect -733 264 -731 269
rect -677 264 -675 269
rect -653 264 -651 269
rect -629 264 -627 269
rect -781 249 -779 254
rect -757 250 -755 255
rect -807 243 -805 248
rect -708 247 -706 257
rect -653 250 -651 255
rect -629 249 -627 254
rect -570 252 -568 257
rect -546 252 -544 257
rect -522 252 -520 257
rect -394 252 -392 257
rect -370 252 -368 257
rect -346 252 -344 257
rect -603 243 -601 248
rect -257 252 -255 257
rect -233 252 -231 257
rect -209 252 -207 257
rect -151 252 -149 257
rect -127 252 -125 257
rect -103 252 -101 257
rect -546 238 -544 243
rect -522 237 -520 242
rect -394 237 -392 242
rect -370 238 -368 243
rect -496 231 -494 236
rect -420 231 -418 236
rect -311 236 -309 246
rect -233 238 -231 243
rect -209 237 -207 242
rect -127 238 -125 243
rect -183 231 -181 236
rect -103 237 -101 242
rect -77 231 -75 236
rect -769 205 -759 207
rect -700 205 -690 207
rect -592 193 -582 195
rect -523 193 -513 195
rect -408 193 -398 195
rect -339 193 -329 195
rect -226 193 -216 195
rect -157 193 -147 195
rect -56 179 -54 184
rect -32 179 -30 184
rect -8 179 -6 184
rect -762 175 -752 177
rect -693 175 -683 177
rect -32 165 -30 170
rect -585 163 -575 165
rect -516 163 -506 165
rect -401 163 -391 165
rect -332 163 -322 165
rect -219 163 -209 165
rect -150 163 -140 165
rect -8 164 -6 169
rect 18 158 20 163
rect -758 131 -756 141
rect -689 131 -687 141
rect -581 119 -579 129
rect -512 119 -510 129
rect -397 119 -395 129
rect -328 119 -326 129
rect -215 119 -213 129
rect -146 119 -144 129
rect -66 101 -64 106
rect -42 101 -40 106
rect -18 101 -16 106
rect -789 46 -787 56
rect -764 47 -762 87
rect -743 47 -741 87
rect -722 47 -720 87
rect -701 47 -699 87
rect -42 87 -40 92
rect -18 86 -16 91
rect 8 80 10 85
rect -665 55 -663 75
rect -635 55 -633 75
rect -488 43 -486 63
rect -458 43 -456 63
rect -304 43 -302 63
rect -274 43 -272 63
rect -122 43 -120 63
rect -92 43 -90 63
rect -489 12 -479 14
rect -236 18 -216 20
rect -17 23 -15 28
rect 7 23 9 28
rect 31 23 33 28
rect -305 12 -295 14
rect 66 18 68 28
rect -123 12 -113 14
rect -17 8 -15 13
rect 7 9 9 14
rect -43 2 -41 7
rect -856 -62 -854 -52
rect -822 -93 -820 -53
rect -801 -93 -799 -53
rect -780 -93 -778 -53
rect -759 -93 -757 -53
rect -694 -64 -692 -44
rect -674 -64 -672 -44
rect -641 -48 -639 -8
rect -620 -48 -618 -8
rect -599 -48 -597 -8
rect -578 -48 -576 -8
rect -419 -30 -417 0
rect -398 -30 -396 0
rect -377 -30 -375 0
rect -236 -2 -216 0
rect -476 -68 -474 -48
rect -456 -68 -454 -48
rect -292 -68 -290 -48
rect -272 -68 -270 -48
rect -110 -68 -108 -48
rect -90 -68 -88 -48
rect -53 -64 -51 -59
rect -29 -64 -27 -59
rect -5 -64 -3 -59
rect -775 -113 -755 -111
rect -29 -78 -27 -73
rect -5 -79 -3 -74
rect -775 -133 -755 -131
rect -731 -170 -729 -130
rect -710 -170 -708 -130
rect -689 -170 -687 -130
rect -668 -170 -666 -130
rect -638 -149 -636 -119
rect -617 -149 -615 -119
rect -596 -149 -594 -119
rect -553 -124 -551 -94
rect -532 -124 -530 -94
rect -511 -124 -509 -94
rect -369 -121 -367 -91
rect -348 -121 -346 -91
rect -327 -121 -325 -91
rect 21 -85 23 -80
rect -190 -117 -188 -112
rect -166 -117 -164 -112
rect -142 -117 -140 -112
rect 21 -112 23 -107
rect -29 -119 -27 -114
rect -5 -118 -3 -113
rect -462 -170 -460 -130
rect -441 -170 -439 -130
rect -420 -170 -418 -130
rect -399 -170 -397 -130
rect -190 -132 -188 -127
rect -166 -131 -164 -126
rect -216 -138 -214 -133
rect -53 -133 -51 -128
rect -29 -133 -27 -128
rect -5 -133 -3 -128
rect -147 -167 -137 -165
rect -630 -177 -610 -175
rect -809 -192 -807 -187
rect -785 -192 -783 -187
rect -761 -192 -759 -187
rect -630 -199 -610 -197
rect -809 -207 -807 -202
rect -785 -206 -783 -201
rect -835 -213 -833 -208
rect -723 -221 -713 -219
<< ptransistor >>
rect -807 284 -805 294
rect -781 284 -779 294
rect -757 284 -755 294
rect -733 283 -731 293
rect -807 260 -805 270
rect -708 272 -706 292
rect -677 283 -675 293
rect -653 284 -651 294
rect -629 284 -627 294
rect -603 284 -601 294
rect -570 271 -568 281
rect -546 272 -544 282
rect -522 272 -520 282
rect -496 272 -494 282
rect -420 272 -418 282
rect -394 272 -392 282
rect -370 272 -368 282
rect -603 260 -601 270
rect -346 271 -344 281
rect -496 248 -494 258
rect -420 248 -418 258
rect -311 261 -309 281
rect -257 271 -255 281
rect -233 272 -231 282
rect -209 272 -207 282
rect -183 272 -181 282
rect -151 271 -149 281
rect -127 272 -125 282
rect -103 272 -101 282
rect -77 272 -75 282
rect -183 248 -181 258
rect -77 248 -75 258
rect -744 205 -724 207
rect -672 205 -652 207
rect -56 198 -54 208
rect -32 199 -30 209
rect -8 199 -6 209
rect 18 199 20 209
rect -567 193 -547 195
rect -495 193 -475 195
rect -383 193 -363 195
rect -311 193 -291 195
rect -201 193 -181 195
rect -129 193 -109 195
rect -737 175 -717 177
rect -665 175 -645 177
rect 18 175 20 185
rect -560 163 -540 165
rect -488 163 -468 165
rect -376 163 -356 165
rect -304 163 -284 165
rect -194 163 -174 165
rect -122 163 -102 165
rect -732 131 -730 151
rect -660 131 -658 151
rect -555 119 -553 139
rect -483 119 -481 139
rect -371 119 -369 139
rect -299 119 -297 139
rect -189 119 -187 139
rect -117 119 -115 139
rect -66 120 -64 130
rect -42 121 -40 131
rect -18 121 -16 131
rect 8 121 10 131
rect -665 89 -663 109
rect -635 89 -633 109
rect 8 97 10 107
rect -488 77 -486 97
rect -458 77 -456 97
rect -304 77 -302 97
rect -274 77 -272 97
rect -122 77 -120 97
rect -92 77 -90 97
rect -43 43 -41 53
rect -17 43 -15 53
rect 7 43 9 53
rect 31 42 33 52
rect 66 43 68 63
rect -789 12 -787 32
rect -764 12 -762 32
rect -743 12 -741 32
rect -722 12 -720 32
rect -701 12 -699 32
rect -641 7 -639 27
rect -620 7 -618 27
rect -599 7 -597 27
rect -578 7 -576 27
rect -419 15 -417 35
rect -398 15 -396 35
rect -377 15 -375 35
rect -464 12 -444 14
rect -202 18 -182 20
rect -43 19 -41 29
rect -280 12 -260 14
rect -98 12 -78 14
rect -856 -37 -854 -17
rect -822 -38 -820 -18
rect -801 -38 -799 -18
rect -780 -38 -778 -18
rect -759 -38 -757 -18
rect -694 -30 -692 -10
rect -674 -30 -672 -10
rect -476 -34 -474 -14
rect -456 -34 -454 -14
rect -202 -2 -182 0
rect -292 -34 -290 -14
rect -272 -34 -270 -14
rect -110 -34 -108 -14
rect -90 -34 -88 -14
rect -53 -45 -51 -35
rect -29 -44 -27 -34
rect -5 -44 -3 -34
rect 21 -44 23 -34
rect -553 -79 -551 -59
rect -532 -79 -530 -59
rect -511 -79 -509 -59
rect -369 -76 -367 -56
rect -348 -76 -346 -56
rect -327 -76 -325 -56
rect 21 -68 23 -58
rect -809 -113 -789 -111
rect -731 -115 -729 -95
rect -710 -115 -708 -95
rect -689 -115 -687 -95
rect -668 -115 -666 -95
rect -638 -104 -636 -84
rect -617 -104 -615 -84
rect -596 -104 -594 -84
rect -809 -133 -789 -131
rect -835 -172 -833 -162
rect -809 -172 -807 -162
rect -785 -172 -783 -162
rect -761 -173 -759 -163
rect -462 -115 -460 -95
rect -441 -115 -439 -95
rect -420 -115 -418 -95
rect -399 -115 -397 -95
rect -216 -97 -214 -87
rect -190 -97 -188 -87
rect -166 -97 -164 -87
rect -142 -98 -140 -88
rect -216 -121 -214 -111
rect 21 -134 23 -124
rect -53 -157 -51 -147
rect -29 -158 -27 -148
rect -5 -158 -3 -148
rect 21 -158 23 -148
rect -122 -167 -102 -165
rect -835 -196 -833 -186
rect -596 -177 -576 -175
rect -596 -199 -576 -197
rect -758 -221 -738 -219
<< ndiffusion >>
rect -782 264 -781 269
rect -779 264 -778 269
rect -758 264 -757 269
rect -755 264 -754 269
rect -734 264 -733 269
rect -731 264 -730 269
rect -678 264 -677 269
rect -675 264 -674 269
rect -654 264 -653 269
rect -651 264 -650 269
rect -630 264 -629 269
rect -627 264 -626 269
rect -782 249 -781 254
rect -779 249 -778 254
rect -758 250 -757 255
rect -755 250 -754 255
rect -808 243 -807 248
rect -805 243 -804 248
rect -709 247 -708 257
rect -706 247 -705 257
rect -654 250 -653 255
rect -651 250 -650 255
rect -630 249 -629 254
rect -627 249 -626 254
rect -571 252 -570 257
rect -568 252 -567 257
rect -547 252 -546 257
rect -544 252 -543 257
rect -523 252 -522 257
rect -520 252 -519 257
rect -395 252 -394 257
rect -392 252 -391 257
rect -371 252 -370 257
rect -368 252 -367 257
rect -347 252 -346 257
rect -344 252 -343 257
rect -604 243 -603 248
rect -601 243 -600 248
rect -258 252 -257 257
rect -255 252 -254 257
rect -234 252 -233 257
rect -231 252 -230 257
rect -210 252 -209 257
rect -207 252 -206 257
rect -152 252 -151 257
rect -149 252 -148 257
rect -128 252 -127 257
rect -125 252 -124 257
rect -104 252 -103 257
rect -101 252 -100 257
rect -547 238 -546 243
rect -544 238 -543 243
rect -523 237 -522 242
rect -520 237 -519 242
rect -395 237 -394 242
rect -392 237 -391 242
rect -371 238 -370 243
rect -368 238 -367 243
rect -497 231 -496 236
rect -494 231 -493 236
rect -421 231 -420 236
rect -418 231 -417 236
rect -312 236 -311 246
rect -309 236 -308 246
rect -234 238 -233 243
rect -231 238 -230 243
rect -210 237 -209 242
rect -207 237 -206 242
rect -128 238 -127 243
rect -125 238 -124 243
rect -184 231 -183 236
rect -181 231 -180 236
rect -104 237 -103 242
rect -101 237 -100 242
rect -78 231 -77 236
rect -75 231 -74 236
rect -769 207 -759 208
rect -700 207 -690 208
rect -769 204 -759 205
rect -700 204 -690 205
rect -592 195 -582 196
rect -523 195 -513 196
rect -408 195 -398 196
rect -339 195 -329 196
rect -226 195 -216 196
rect -157 195 -147 196
rect -592 192 -582 193
rect -523 192 -513 193
rect -408 192 -398 193
rect -339 192 -329 193
rect -226 192 -216 193
rect -157 192 -147 193
rect -762 177 -752 178
rect -693 177 -683 178
rect -57 179 -56 184
rect -54 179 -53 184
rect -33 179 -32 184
rect -30 179 -29 184
rect -9 179 -8 184
rect -6 179 -5 184
rect -762 174 -752 175
rect -693 174 -683 175
rect -585 165 -575 166
rect -516 165 -506 166
rect -401 165 -391 166
rect -332 165 -322 166
rect -219 165 -209 166
rect -150 165 -140 166
rect -33 165 -32 170
rect -30 165 -29 170
rect -585 162 -575 163
rect -516 162 -506 163
rect -401 162 -391 163
rect -332 162 -322 163
rect -219 162 -209 163
rect -150 162 -140 163
rect -9 164 -8 169
rect -6 164 -5 169
rect 17 158 18 163
rect 20 158 21 163
rect -759 131 -758 141
rect -756 131 -755 141
rect -690 131 -689 141
rect -687 131 -686 141
rect -582 119 -581 129
rect -579 119 -578 129
rect -513 119 -512 129
rect -510 119 -509 129
rect -398 119 -397 129
rect -395 119 -394 129
rect -329 119 -328 129
rect -326 119 -325 129
rect -216 119 -215 129
rect -213 119 -212 129
rect -147 119 -146 129
rect -144 119 -143 129
rect -67 101 -66 106
rect -64 101 -63 106
rect -43 101 -42 106
rect -40 101 -39 106
rect -19 101 -18 106
rect -16 101 -15 106
rect -790 46 -789 56
rect -787 46 -786 56
rect -765 47 -764 87
rect -762 47 -761 87
rect -744 47 -743 87
rect -741 47 -740 87
rect -723 47 -722 87
rect -720 47 -719 87
rect -702 47 -701 87
rect -699 47 -698 87
rect -43 87 -42 92
rect -40 87 -39 92
rect -19 86 -18 91
rect -16 86 -15 91
rect 7 80 8 85
rect 10 80 11 85
rect -666 55 -665 75
rect -663 55 -662 75
rect -636 55 -635 75
rect -633 55 -632 75
rect -489 43 -488 63
rect -486 43 -485 63
rect -459 43 -458 63
rect -456 43 -455 63
rect -305 43 -304 63
rect -302 43 -301 63
rect -275 43 -274 63
rect -272 43 -271 63
rect -123 43 -122 63
rect -120 43 -119 63
rect -93 43 -92 63
rect -90 43 -89 63
rect -489 14 -479 15
rect -236 20 -216 21
rect -489 11 -479 12
rect -305 14 -295 15
rect -18 23 -17 28
rect -15 23 -14 28
rect 6 23 7 28
rect 9 23 10 28
rect 30 23 31 28
rect 33 23 34 28
rect -236 17 -216 18
rect -123 14 -113 15
rect 65 18 66 28
rect 68 18 69 28
rect -305 11 -295 12
rect -123 11 -113 12
rect -18 8 -17 13
rect -15 8 -14 13
rect 6 9 7 14
rect 9 9 10 14
rect -236 0 -216 1
rect -44 2 -43 7
rect -41 2 -40 7
rect -857 -62 -856 -52
rect -854 -62 -853 -52
rect -823 -93 -822 -53
rect -820 -93 -819 -53
rect -802 -93 -801 -53
rect -799 -93 -798 -53
rect -781 -93 -780 -53
rect -778 -93 -777 -53
rect -760 -93 -759 -53
rect -757 -93 -756 -53
rect -695 -64 -694 -44
rect -692 -64 -691 -44
rect -675 -64 -674 -44
rect -672 -64 -671 -44
rect -642 -48 -641 -8
rect -639 -48 -638 -8
rect -621 -48 -620 -8
rect -618 -48 -617 -8
rect -600 -48 -599 -8
rect -597 -48 -596 -8
rect -579 -48 -578 -8
rect -576 -48 -575 -8
rect -420 -30 -419 0
rect -417 -30 -416 0
rect -399 -30 -398 0
rect -396 -30 -395 0
rect -378 -30 -377 0
rect -375 -30 -374 0
rect -236 -3 -216 -2
rect -477 -68 -476 -48
rect -474 -68 -473 -48
rect -457 -68 -456 -48
rect -454 -68 -453 -48
rect -293 -68 -292 -48
rect -290 -68 -289 -48
rect -273 -68 -272 -48
rect -270 -68 -269 -48
rect -111 -68 -110 -48
rect -108 -68 -107 -48
rect -91 -68 -90 -48
rect -88 -68 -87 -48
rect -54 -64 -53 -59
rect -51 -64 -50 -59
rect -30 -64 -29 -59
rect -27 -64 -26 -59
rect -6 -64 -5 -59
rect -3 -64 -2 -59
rect -775 -111 -755 -110
rect -775 -114 -755 -113
rect -30 -78 -29 -73
rect -27 -78 -26 -73
rect -6 -79 -5 -74
rect -3 -79 -2 -74
rect -775 -131 -755 -130
rect -775 -134 -755 -133
rect -732 -170 -731 -130
rect -729 -170 -728 -130
rect -711 -170 -710 -130
rect -708 -170 -707 -130
rect -690 -170 -689 -130
rect -687 -170 -686 -130
rect -669 -170 -668 -130
rect -666 -170 -665 -130
rect -639 -149 -638 -119
rect -636 -149 -635 -119
rect -618 -149 -617 -119
rect -615 -149 -614 -119
rect -597 -149 -596 -119
rect -594 -149 -593 -119
rect -554 -124 -553 -94
rect -551 -124 -550 -94
rect -533 -124 -532 -94
rect -530 -124 -529 -94
rect -512 -124 -511 -94
rect -509 -124 -508 -94
rect -370 -121 -369 -91
rect -367 -121 -366 -91
rect -349 -121 -348 -91
rect -346 -121 -345 -91
rect -328 -121 -327 -91
rect -325 -121 -324 -91
rect 20 -85 21 -80
rect 23 -85 24 -80
rect -191 -117 -190 -112
rect -188 -117 -187 -112
rect -167 -117 -166 -112
rect -164 -117 -163 -112
rect -143 -117 -142 -112
rect -140 -117 -139 -112
rect 20 -112 21 -107
rect 23 -112 24 -107
rect -30 -119 -29 -114
rect -27 -119 -26 -114
rect -6 -118 -5 -113
rect -3 -118 -2 -113
rect -463 -170 -462 -130
rect -460 -170 -459 -130
rect -442 -170 -441 -130
rect -439 -170 -438 -130
rect -421 -170 -420 -130
rect -418 -170 -417 -130
rect -400 -170 -399 -130
rect -397 -170 -396 -130
rect -191 -132 -190 -127
rect -188 -132 -187 -127
rect -167 -131 -166 -126
rect -164 -131 -163 -126
rect -217 -138 -216 -133
rect -214 -138 -213 -133
rect -54 -133 -53 -128
rect -51 -133 -50 -128
rect -30 -133 -29 -128
rect -27 -133 -26 -128
rect -6 -133 -5 -128
rect -3 -133 -2 -128
rect -147 -165 -137 -164
rect -147 -168 -137 -167
rect -630 -175 -610 -174
rect -630 -178 -610 -177
rect -810 -192 -809 -187
rect -807 -192 -806 -187
rect -786 -192 -785 -187
rect -783 -192 -782 -187
rect -762 -192 -761 -187
rect -759 -192 -758 -187
rect -630 -197 -610 -196
rect -630 -200 -610 -199
rect -810 -207 -809 -202
rect -807 -207 -806 -202
rect -786 -206 -785 -201
rect -783 -206 -782 -201
rect -836 -213 -835 -208
rect -833 -213 -832 -208
rect -723 -219 -713 -218
rect -723 -222 -713 -221
<< pdiffusion >>
rect -808 284 -807 294
rect -805 284 -804 294
rect -782 284 -781 294
rect -779 284 -778 294
rect -758 284 -757 294
rect -755 284 -754 294
rect -734 283 -733 293
rect -731 283 -730 293
rect -808 260 -807 270
rect -805 260 -804 270
rect -709 272 -708 292
rect -706 272 -705 292
rect -678 283 -677 293
rect -675 283 -674 293
rect -654 284 -653 294
rect -651 284 -650 294
rect -630 284 -629 294
rect -627 284 -626 294
rect -604 284 -603 294
rect -601 284 -600 294
rect -571 271 -570 281
rect -568 271 -567 281
rect -547 272 -546 282
rect -544 272 -543 282
rect -523 272 -522 282
rect -520 272 -519 282
rect -497 272 -496 282
rect -494 272 -493 282
rect -421 272 -420 282
rect -418 272 -417 282
rect -395 272 -394 282
rect -392 272 -391 282
rect -371 272 -370 282
rect -368 272 -367 282
rect -604 260 -603 270
rect -601 260 -600 270
rect -347 271 -346 281
rect -344 271 -343 281
rect -497 248 -496 258
rect -494 248 -493 258
rect -421 248 -420 258
rect -418 248 -417 258
rect -312 261 -311 281
rect -309 261 -308 281
rect -258 271 -257 281
rect -255 271 -254 281
rect -234 272 -233 282
rect -231 272 -230 282
rect -210 272 -209 282
rect -207 272 -206 282
rect -184 272 -183 282
rect -181 272 -180 282
rect -152 271 -151 281
rect -149 271 -148 281
rect -128 272 -127 282
rect -125 272 -124 282
rect -104 272 -103 282
rect -101 272 -100 282
rect -78 272 -77 282
rect -75 272 -74 282
rect -184 248 -183 258
rect -181 248 -180 258
rect -78 248 -77 258
rect -75 248 -74 258
rect -744 207 -724 208
rect -672 207 -652 208
rect -744 204 -724 205
rect -672 204 -652 205
rect -567 195 -547 196
rect -495 195 -475 196
rect -383 195 -363 196
rect -311 195 -291 196
rect -201 195 -181 196
rect -57 198 -56 208
rect -54 198 -53 208
rect -33 199 -32 209
rect -30 199 -29 209
rect -9 199 -8 209
rect -6 199 -5 209
rect 17 199 18 209
rect 20 199 21 209
rect -129 195 -109 196
rect -567 192 -547 193
rect -495 192 -475 193
rect -383 192 -363 193
rect -311 192 -291 193
rect -201 192 -181 193
rect -129 192 -109 193
rect -737 177 -717 178
rect -665 177 -645 178
rect 17 175 18 185
rect 20 175 21 185
rect -737 174 -717 175
rect -665 174 -645 175
rect -560 165 -540 166
rect -488 165 -468 166
rect -376 165 -356 166
rect -304 165 -284 166
rect -194 165 -174 166
rect -122 165 -102 166
rect -560 162 -540 163
rect -488 162 -468 163
rect -376 162 -356 163
rect -304 162 -284 163
rect -194 162 -174 163
rect -122 162 -102 163
rect -733 131 -732 151
rect -730 131 -729 151
rect -661 131 -660 151
rect -658 131 -657 151
rect -556 119 -555 139
rect -553 119 -552 139
rect -484 119 -483 139
rect -481 119 -480 139
rect -372 119 -371 139
rect -369 119 -368 139
rect -300 119 -299 139
rect -297 119 -296 139
rect -190 119 -189 139
rect -187 119 -186 139
rect -118 119 -117 139
rect -115 119 -114 139
rect -67 120 -66 130
rect -64 120 -63 130
rect -43 121 -42 131
rect -40 121 -39 131
rect -19 121 -18 131
rect -16 121 -15 131
rect 7 121 8 131
rect 10 121 11 131
rect -666 89 -665 109
rect -663 89 -662 109
rect -636 89 -635 109
rect -633 89 -632 109
rect 7 97 8 107
rect 10 97 11 107
rect -489 77 -488 97
rect -486 77 -485 97
rect -459 77 -458 97
rect -456 77 -455 97
rect -305 77 -304 97
rect -302 77 -301 97
rect -275 77 -274 97
rect -272 77 -271 97
rect -123 77 -122 97
rect -120 77 -119 97
rect -93 77 -92 97
rect -90 77 -89 97
rect -44 43 -43 53
rect -41 43 -40 53
rect -18 43 -17 53
rect -15 43 -14 53
rect 6 43 7 53
rect 9 43 10 53
rect 30 42 31 52
rect 33 42 34 52
rect 65 43 66 63
rect 68 43 69 63
rect -790 12 -789 32
rect -787 12 -786 32
rect -765 12 -764 32
rect -762 12 -761 32
rect -744 12 -743 32
rect -741 12 -740 32
rect -723 12 -722 32
rect -720 12 -719 32
rect -702 12 -701 32
rect -699 12 -698 32
rect -642 7 -641 27
rect -639 7 -638 27
rect -621 7 -620 27
rect -618 7 -617 27
rect -600 7 -599 27
rect -597 7 -596 27
rect -579 7 -578 27
rect -576 7 -575 27
rect -420 15 -419 35
rect -417 15 -416 35
rect -399 15 -398 35
rect -396 15 -395 35
rect -378 15 -377 35
rect -375 15 -374 35
rect -202 20 -182 21
rect -464 14 -444 15
rect -464 11 -444 12
rect -44 19 -43 29
rect -41 19 -40 29
rect -280 14 -260 15
rect -202 17 -182 18
rect -98 14 -78 15
rect -280 11 -260 12
rect -98 11 -78 12
rect -202 0 -182 1
rect -857 -37 -856 -17
rect -854 -37 -853 -17
rect -823 -38 -822 -18
rect -820 -38 -819 -18
rect -802 -38 -801 -18
rect -799 -38 -798 -18
rect -781 -38 -780 -18
rect -778 -38 -777 -18
rect -760 -38 -759 -18
rect -757 -38 -756 -18
rect -695 -30 -694 -10
rect -692 -30 -691 -10
rect -675 -30 -674 -10
rect -672 -30 -671 -10
rect -477 -34 -476 -14
rect -474 -34 -473 -14
rect -457 -34 -456 -14
rect -454 -34 -453 -14
rect -202 -3 -182 -2
rect -293 -34 -292 -14
rect -290 -34 -289 -14
rect -273 -34 -272 -14
rect -270 -34 -269 -14
rect -111 -34 -110 -14
rect -108 -34 -107 -14
rect -91 -34 -90 -14
rect -88 -34 -87 -14
rect -54 -45 -53 -35
rect -51 -45 -50 -35
rect -30 -44 -29 -34
rect -27 -44 -26 -34
rect -6 -44 -5 -34
rect -3 -44 -2 -34
rect 20 -44 21 -34
rect 23 -44 24 -34
rect -554 -79 -553 -59
rect -551 -79 -550 -59
rect -533 -79 -532 -59
rect -530 -79 -529 -59
rect -512 -79 -511 -59
rect -509 -79 -508 -59
rect -370 -76 -369 -56
rect -367 -76 -366 -56
rect -349 -76 -348 -56
rect -346 -76 -345 -56
rect -328 -76 -327 -56
rect -325 -76 -324 -56
rect 20 -68 21 -58
rect 23 -68 24 -58
rect -809 -111 -789 -110
rect -809 -114 -789 -113
rect -732 -115 -731 -95
rect -729 -115 -728 -95
rect -711 -115 -710 -95
rect -708 -115 -707 -95
rect -690 -115 -689 -95
rect -687 -115 -686 -95
rect -669 -115 -668 -95
rect -666 -115 -665 -95
rect -639 -104 -638 -84
rect -636 -104 -635 -84
rect -618 -104 -617 -84
rect -615 -104 -614 -84
rect -597 -104 -596 -84
rect -594 -104 -593 -84
rect -809 -131 -789 -130
rect -809 -134 -789 -133
rect -836 -172 -835 -162
rect -833 -172 -832 -162
rect -810 -172 -809 -162
rect -807 -172 -806 -162
rect -786 -172 -785 -162
rect -783 -172 -782 -162
rect -762 -173 -761 -163
rect -759 -173 -758 -163
rect -463 -115 -462 -95
rect -460 -115 -459 -95
rect -442 -115 -441 -95
rect -439 -115 -438 -95
rect -421 -115 -420 -95
rect -418 -115 -417 -95
rect -400 -115 -399 -95
rect -397 -115 -396 -95
rect -217 -97 -216 -87
rect -214 -97 -213 -87
rect -191 -97 -190 -87
rect -188 -97 -187 -87
rect -167 -97 -166 -87
rect -164 -97 -163 -87
rect -143 -98 -142 -88
rect -140 -98 -139 -88
rect -217 -121 -216 -111
rect -214 -121 -213 -111
rect 20 -134 21 -124
rect 23 -134 24 -124
rect -54 -157 -53 -147
rect -51 -157 -50 -147
rect -30 -158 -29 -148
rect -27 -158 -26 -148
rect -6 -158 -5 -148
rect -3 -158 -2 -148
rect 20 -158 21 -148
rect 23 -158 24 -148
rect -122 -165 -102 -164
rect -836 -196 -835 -186
rect -833 -196 -832 -186
rect -122 -168 -102 -167
rect -596 -175 -576 -174
rect -596 -178 -576 -177
rect -596 -197 -576 -196
rect -596 -200 -576 -199
rect -758 -219 -738 -218
rect -758 -222 -738 -221
<< ndcontact >>
rect -786 264 -782 269
rect -778 264 -774 269
rect -762 264 -758 269
rect -754 264 -750 269
rect -738 264 -734 269
rect -730 264 -726 269
rect -682 264 -678 269
rect -674 264 -670 269
rect -658 264 -654 269
rect -650 264 -646 269
rect -634 264 -630 269
rect -626 264 -622 269
rect -786 249 -782 254
rect -778 249 -774 254
rect -762 250 -758 255
rect -754 250 -750 255
rect -812 243 -808 248
rect -804 243 -800 248
rect -713 247 -709 257
rect -705 247 -701 257
rect -658 250 -654 255
rect -650 250 -646 255
rect -634 249 -630 254
rect -626 249 -622 254
rect -575 252 -571 257
rect -567 252 -563 257
rect -551 252 -547 257
rect -543 252 -539 257
rect -527 252 -523 257
rect -519 252 -515 257
rect -399 252 -395 257
rect -391 252 -387 257
rect -375 252 -371 257
rect -367 252 -363 257
rect -351 252 -347 257
rect -343 252 -339 257
rect -608 243 -604 248
rect -600 243 -596 248
rect -262 252 -258 257
rect -254 252 -250 257
rect -238 252 -234 257
rect -230 252 -226 257
rect -214 252 -210 257
rect -206 252 -202 257
rect -156 252 -152 257
rect -148 252 -144 257
rect -132 252 -128 257
rect -124 252 -120 257
rect -108 252 -104 257
rect -100 252 -96 257
rect -551 238 -547 243
rect -543 238 -539 243
rect -527 237 -523 242
rect -519 237 -515 242
rect -399 237 -395 242
rect -391 237 -387 242
rect -375 238 -371 243
rect -367 238 -363 243
rect -501 231 -497 236
rect -493 231 -489 236
rect -425 231 -421 236
rect -417 231 -413 236
rect -316 236 -312 246
rect -308 236 -304 246
rect -238 238 -234 243
rect -230 238 -226 243
rect -214 237 -210 242
rect -206 237 -202 242
rect -132 238 -128 243
rect -124 238 -120 243
rect -188 231 -184 236
rect -180 231 -176 236
rect -108 237 -104 242
rect -100 237 -96 242
rect -82 231 -78 236
rect -74 231 -70 236
rect -769 208 -759 212
rect -700 208 -690 212
rect -769 200 -759 204
rect -700 200 -690 204
rect -592 196 -582 200
rect -523 196 -513 200
rect -408 196 -398 200
rect -339 196 -329 200
rect -226 196 -216 200
rect -157 196 -147 200
rect -592 188 -582 192
rect -523 188 -513 192
rect -408 188 -398 192
rect -339 188 -329 192
rect -226 188 -216 192
rect -157 188 -147 192
rect -762 178 -752 182
rect -693 178 -683 182
rect -61 179 -57 184
rect -53 179 -49 184
rect -37 179 -33 184
rect -29 179 -25 184
rect -13 179 -9 184
rect -5 179 -1 184
rect -762 170 -752 174
rect -693 170 -683 174
rect -585 166 -575 170
rect -516 166 -506 170
rect -401 166 -391 170
rect -332 166 -322 170
rect -219 166 -209 170
rect -150 166 -140 170
rect -37 165 -33 170
rect -29 165 -25 170
rect -585 158 -575 162
rect -516 158 -506 162
rect -401 158 -391 162
rect -332 158 -322 162
rect -219 158 -209 162
rect -150 158 -140 162
rect -13 164 -9 169
rect -5 164 -1 169
rect 13 158 17 163
rect 21 158 25 163
rect -763 131 -759 141
rect -755 131 -751 141
rect -694 131 -690 141
rect -686 131 -682 141
rect -586 119 -582 129
rect -578 119 -574 129
rect -517 119 -513 129
rect -509 119 -505 129
rect -402 119 -398 129
rect -394 119 -390 129
rect -333 119 -329 129
rect -325 119 -321 129
rect -220 119 -216 129
rect -212 119 -208 129
rect -151 119 -147 129
rect -143 119 -139 129
rect -71 101 -67 106
rect -63 101 -59 106
rect -47 101 -43 106
rect -39 101 -35 106
rect -23 101 -19 106
rect -15 101 -11 106
rect -794 46 -790 56
rect -786 46 -782 56
rect -769 47 -765 87
rect -761 47 -757 87
rect -748 47 -744 87
rect -740 47 -736 87
rect -727 47 -723 87
rect -719 47 -715 87
rect -706 47 -702 87
rect -698 47 -694 87
rect -47 87 -43 92
rect -39 87 -35 92
rect -23 86 -19 91
rect -15 86 -11 91
rect 3 80 7 85
rect 11 80 15 85
rect -670 55 -666 75
rect -662 55 -658 75
rect -640 55 -636 75
rect -632 55 -628 75
rect -493 43 -489 63
rect -485 43 -481 63
rect -463 43 -459 63
rect -455 43 -451 63
rect -309 43 -305 63
rect -301 43 -297 63
rect -279 43 -275 63
rect -271 43 -267 63
rect -127 43 -123 63
rect -119 43 -115 63
rect -97 43 -93 63
rect -89 43 -85 63
rect -489 15 -479 19
rect -236 21 -216 25
rect -305 15 -295 19
rect -489 7 -479 11
rect -22 23 -18 28
rect -14 23 -10 28
rect 2 23 6 28
rect 10 23 14 28
rect 26 23 30 28
rect 34 23 38 28
rect -236 13 -216 17
rect -123 15 -113 19
rect 61 18 65 28
rect 69 18 73 28
rect -305 7 -295 11
rect -123 7 -113 11
rect -22 8 -18 13
rect -14 8 -10 13
rect 2 9 6 14
rect 10 9 14 14
rect -236 1 -216 5
rect -48 2 -44 7
rect -40 2 -36 7
rect -861 -62 -857 -52
rect -853 -62 -849 -52
rect -827 -93 -823 -53
rect -819 -93 -815 -53
rect -806 -93 -802 -53
rect -798 -93 -794 -53
rect -785 -93 -781 -53
rect -777 -93 -773 -53
rect -764 -93 -760 -53
rect -756 -93 -752 -53
rect -699 -64 -695 -44
rect -691 -64 -687 -44
rect -679 -64 -675 -44
rect -671 -64 -667 -44
rect -646 -48 -642 -8
rect -638 -48 -634 -8
rect -625 -48 -621 -8
rect -617 -48 -613 -8
rect -604 -48 -600 -8
rect -596 -48 -592 -8
rect -583 -48 -579 -8
rect -575 -48 -571 -8
rect -424 -30 -420 0
rect -416 -30 -412 0
rect -403 -30 -399 0
rect -395 -30 -391 0
rect -382 -30 -378 0
rect -374 -30 -370 0
rect -236 -7 -216 -3
rect -481 -68 -477 -48
rect -473 -68 -469 -48
rect -461 -68 -457 -48
rect -453 -68 -449 -48
rect -297 -68 -293 -48
rect -289 -68 -285 -48
rect -277 -68 -273 -48
rect -269 -68 -265 -48
rect -115 -68 -111 -48
rect -107 -68 -103 -48
rect -95 -68 -91 -48
rect -87 -68 -83 -48
rect -58 -64 -54 -59
rect -50 -64 -46 -59
rect -34 -64 -30 -59
rect -26 -64 -22 -59
rect -10 -64 -6 -59
rect -2 -64 2 -59
rect -775 -110 -755 -106
rect -775 -118 -755 -114
rect -34 -78 -30 -73
rect -26 -78 -22 -73
rect -10 -79 -6 -74
rect -2 -79 2 -74
rect -775 -130 -755 -126
rect -775 -138 -755 -134
rect -736 -170 -732 -130
rect -728 -170 -724 -130
rect -715 -170 -711 -130
rect -707 -170 -703 -130
rect -694 -170 -690 -130
rect -686 -170 -682 -130
rect -673 -170 -669 -130
rect -665 -170 -661 -130
rect -643 -149 -639 -119
rect -635 -149 -631 -119
rect -622 -149 -618 -119
rect -614 -149 -610 -119
rect -601 -149 -597 -119
rect -593 -149 -589 -119
rect -558 -124 -554 -94
rect -550 -124 -546 -94
rect -537 -124 -533 -94
rect -529 -124 -525 -94
rect -516 -124 -512 -94
rect -508 -124 -504 -94
rect -374 -121 -370 -91
rect -366 -121 -362 -91
rect -353 -121 -349 -91
rect -345 -121 -341 -91
rect -332 -121 -328 -91
rect -324 -121 -320 -91
rect 16 -85 20 -80
rect 24 -85 28 -80
rect -195 -117 -191 -112
rect -187 -117 -183 -112
rect -171 -117 -167 -112
rect -163 -117 -159 -112
rect -147 -117 -143 -112
rect -139 -117 -135 -112
rect 16 -112 20 -107
rect 24 -112 28 -107
rect -34 -119 -30 -114
rect -26 -119 -22 -114
rect -10 -118 -6 -113
rect -2 -118 2 -113
rect -467 -170 -463 -130
rect -459 -170 -455 -130
rect -446 -170 -442 -130
rect -438 -170 -434 -130
rect -425 -170 -421 -130
rect -417 -170 -413 -130
rect -404 -170 -400 -130
rect -396 -170 -392 -130
rect -195 -132 -191 -127
rect -187 -132 -183 -127
rect -171 -131 -167 -126
rect -163 -131 -159 -126
rect -221 -138 -217 -133
rect -213 -138 -209 -133
rect -58 -133 -54 -128
rect -50 -133 -46 -128
rect -34 -133 -30 -128
rect -26 -133 -22 -128
rect -10 -133 -6 -128
rect -2 -133 2 -128
rect -147 -164 -137 -160
rect -630 -174 -610 -170
rect -147 -172 -137 -168
rect -630 -182 -610 -178
rect -814 -192 -810 -187
rect -806 -192 -802 -187
rect -790 -192 -786 -187
rect -782 -192 -778 -187
rect -766 -192 -762 -187
rect -758 -192 -754 -187
rect -630 -196 -610 -192
rect -814 -207 -810 -202
rect -806 -207 -802 -202
rect -790 -206 -786 -201
rect -782 -206 -778 -201
rect -630 -204 -610 -200
rect -840 -213 -836 -208
rect -832 -213 -828 -208
rect -723 -218 -713 -214
rect -723 -226 -713 -222
<< pdcontact >>
rect -812 284 -808 294
rect -804 284 -800 294
rect -786 284 -782 294
rect -778 284 -774 294
rect -762 284 -758 294
rect -754 284 -750 294
rect -738 283 -734 293
rect -730 283 -726 293
rect -812 260 -808 270
rect -804 260 -800 270
rect -713 272 -709 292
rect -705 272 -701 292
rect -682 283 -678 293
rect -674 283 -670 293
rect -658 284 -654 294
rect -650 284 -646 294
rect -634 284 -630 294
rect -626 284 -622 294
rect -608 284 -604 294
rect -600 284 -596 294
rect -575 271 -571 281
rect -567 271 -563 281
rect -551 272 -547 282
rect -543 272 -539 282
rect -527 272 -523 282
rect -519 272 -515 282
rect -501 272 -497 282
rect -493 272 -489 282
rect -425 272 -421 282
rect -417 272 -413 282
rect -399 272 -395 282
rect -391 272 -387 282
rect -375 272 -371 282
rect -367 272 -363 282
rect -608 260 -604 270
rect -600 260 -596 270
rect -351 271 -347 281
rect -343 271 -339 281
rect -501 248 -497 258
rect -493 248 -489 258
rect -425 248 -421 258
rect -417 248 -413 258
rect -316 261 -312 281
rect -308 261 -304 281
rect -262 271 -258 281
rect -254 271 -250 281
rect -238 272 -234 282
rect -230 272 -226 282
rect -214 272 -210 282
rect -206 272 -202 282
rect -188 272 -184 282
rect -180 272 -176 282
rect -156 271 -152 281
rect -148 271 -144 281
rect -132 272 -128 282
rect -124 272 -120 282
rect -108 272 -104 282
rect -100 272 -96 282
rect -82 272 -78 282
rect -74 272 -70 282
rect -188 248 -184 258
rect -180 248 -176 258
rect -82 248 -78 258
rect -74 248 -70 258
rect -744 208 -724 212
rect -672 208 -652 212
rect -744 200 -724 204
rect -672 200 -652 204
rect -567 196 -547 200
rect -495 196 -475 200
rect -383 196 -363 200
rect -311 196 -291 200
rect -201 196 -181 200
rect -129 196 -109 200
rect -61 198 -57 208
rect -53 198 -49 208
rect -37 199 -33 209
rect -29 199 -25 209
rect -13 199 -9 209
rect -5 199 -1 209
rect 13 199 17 209
rect 21 199 25 209
rect -567 188 -547 192
rect -495 188 -475 192
rect -383 188 -363 192
rect -311 188 -291 192
rect -201 188 -181 192
rect -129 188 -109 192
rect -737 178 -717 182
rect -665 178 -645 182
rect 13 175 17 185
rect 21 175 25 185
rect -737 170 -717 174
rect -665 170 -645 174
rect -560 166 -540 170
rect -488 166 -468 170
rect -376 166 -356 170
rect -304 166 -284 170
rect -194 166 -174 170
rect -122 166 -102 170
rect -560 158 -540 162
rect -488 158 -468 162
rect -376 158 -356 162
rect -304 158 -284 162
rect -194 158 -174 162
rect -122 158 -102 162
rect -737 131 -733 151
rect -729 131 -725 151
rect -665 131 -661 151
rect -657 131 -653 151
rect -560 119 -556 139
rect -552 119 -548 139
rect -488 119 -484 139
rect -480 119 -476 139
rect -376 119 -372 139
rect -368 119 -364 139
rect -304 119 -300 139
rect -296 119 -292 139
rect -194 119 -190 139
rect -186 119 -182 139
rect -122 119 -118 139
rect -114 119 -110 139
rect -71 120 -67 130
rect -63 120 -59 130
rect -47 121 -43 131
rect -39 121 -35 131
rect -23 121 -19 131
rect -15 121 -11 131
rect 3 121 7 131
rect 11 121 15 131
rect -670 89 -666 109
rect -662 89 -658 109
rect -640 89 -636 109
rect -632 89 -628 109
rect 3 97 7 107
rect 11 97 15 107
rect -493 77 -489 97
rect -485 77 -481 97
rect -463 77 -459 97
rect -455 77 -451 97
rect -309 77 -305 97
rect -301 77 -297 97
rect -279 77 -275 97
rect -271 77 -267 97
rect -127 77 -123 97
rect -119 77 -115 97
rect -97 77 -93 97
rect -89 77 -85 97
rect -48 43 -44 53
rect -40 43 -36 53
rect -22 43 -18 53
rect -14 43 -10 53
rect 2 43 6 53
rect 10 43 14 53
rect 26 42 30 52
rect 34 42 38 52
rect 61 43 65 63
rect 69 43 73 63
rect -794 12 -790 32
rect -786 12 -782 32
rect -769 12 -765 32
rect -761 12 -757 32
rect -748 12 -744 32
rect -740 12 -736 32
rect -727 12 -723 32
rect -719 12 -715 32
rect -706 12 -702 32
rect -698 12 -694 32
rect -646 7 -642 27
rect -638 7 -634 27
rect -625 7 -621 27
rect -617 7 -613 27
rect -604 7 -600 27
rect -596 7 -592 27
rect -583 7 -579 27
rect -575 7 -571 27
rect -464 15 -444 19
rect -424 15 -420 35
rect -416 15 -412 35
rect -403 15 -399 35
rect -395 15 -391 35
rect -382 15 -378 35
rect -374 15 -370 35
rect -202 21 -182 25
rect -464 7 -444 11
rect -280 15 -260 19
rect -48 19 -44 29
rect -40 19 -36 29
rect -202 13 -182 17
rect -98 15 -78 19
rect -280 7 -260 11
rect -98 7 -78 11
rect -202 1 -182 5
rect -861 -37 -857 -17
rect -853 -37 -849 -17
rect -827 -38 -823 -18
rect -819 -38 -815 -18
rect -806 -38 -802 -18
rect -798 -38 -794 -18
rect -785 -38 -781 -18
rect -777 -38 -773 -18
rect -764 -38 -760 -18
rect -756 -38 -752 -18
rect -699 -30 -695 -10
rect -691 -30 -687 -10
rect -679 -30 -675 -10
rect -671 -30 -667 -10
rect -481 -34 -477 -14
rect -473 -34 -469 -14
rect -461 -34 -457 -14
rect -453 -34 -449 -14
rect -202 -7 -182 -3
rect -297 -34 -293 -14
rect -289 -34 -285 -14
rect -277 -34 -273 -14
rect -269 -34 -265 -14
rect -115 -34 -111 -14
rect -107 -34 -103 -14
rect -95 -34 -91 -14
rect -87 -34 -83 -14
rect -58 -45 -54 -35
rect -50 -45 -46 -35
rect -34 -44 -30 -34
rect -26 -44 -22 -34
rect -10 -44 -6 -34
rect -2 -44 2 -34
rect 16 -44 20 -34
rect 24 -44 28 -34
rect -558 -79 -554 -59
rect -550 -79 -546 -59
rect -537 -79 -533 -59
rect -529 -79 -525 -59
rect -516 -79 -512 -59
rect -508 -79 -504 -59
rect -374 -76 -370 -56
rect -366 -76 -362 -56
rect -353 -76 -349 -56
rect -345 -76 -341 -56
rect -332 -76 -328 -56
rect -324 -76 -320 -56
rect 16 -68 20 -58
rect 24 -68 28 -58
rect -809 -110 -789 -106
rect -809 -118 -789 -114
rect -736 -115 -732 -95
rect -728 -115 -724 -95
rect -715 -115 -711 -95
rect -707 -115 -703 -95
rect -694 -115 -690 -95
rect -686 -115 -682 -95
rect -673 -115 -669 -95
rect -665 -115 -661 -95
rect -643 -104 -639 -84
rect -635 -104 -631 -84
rect -622 -104 -618 -84
rect -614 -104 -610 -84
rect -601 -104 -597 -84
rect -593 -104 -589 -84
rect -809 -130 -789 -126
rect -809 -138 -789 -134
rect -840 -172 -836 -162
rect -832 -172 -828 -162
rect -814 -172 -810 -162
rect -806 -172 -802 -162
rect -790 -172 -786 -162
rect -782 -172 -778 -162
rect -766 -173 -762 -163
rect -758 -173 -754 -163
rect -467 -115 -463 -95
rect -459 -115 -455 -95
rect -446 -115 -442 -95
rect -438 -115 -434 -95
rect -425 -115 -421 -95
rect -417 -115 -413 -95
rect -404 -115 -400 -95
rect -396 -115 -392 -95
rect -221 -97 -217 -87
rect -213 -97 -209 -87
rect -195 -97 -191 -87
rect -187 -97 -183 -87
rect -171 -97 -167 -87
rect -163 -97 -159 -87
rect -147 -98 -143 -88
rect -139 -98 -135 -88
rect -221 -121 -217 -111
rect -213 -121 -209 -111
rect 16 -134 20 -124
rect 24 -134 28 -124
rect -58 -157 -54 -147
rect -50 -157 -46 -147
rect -34 -158 -30 -148
rect -26 -158 -22 -148
rect -10 -158 -6 -148
rect -2 -158 2 -148
rect 16 -158 20 -148
rect 24 -158 28 -148
rect -122 -164 -102 -160
rect -840 -196 -836 -186
rect -832 -196 -828 -186
rect -596 -174 -576 -170
rect -122 -172 -102 -168
rect -596 -182 -576 -178
rect -596 -196 -576 -192
rect -596 -204 -576 -200
rect -758 -218 -738 -214
rect -758 -226 -738 -222
<< polysilicon >>
rect -807 294 -805 297
rect -781 294 -779 297
rect -757 294 -755 297
rect -733 293 -731 296
rect -807 281 -805 284
rect -781 281 -779 284
rect -757 281 -755 284
rect -708 292 -706 295
rect -677 293 -675 296
rect -653 294 -651 297
rect -629 294 -627 297
rect -603 294 -601 297
rect -807 270 -805 273
rect -781 269 -779 272
rect -757 269 -755 272
rect -733 269 -731 283
rect -781 261 -779 264
rect -757 261 -755 264
rect -733 261 -731 264
rect -807 257 -805 260
rect -781 254 -779 257
rect -757 255 -755 258
rect -708 257 -706 272
rect -677 269 -675 283
rect -653 281 -651 284
rect -629 281 -627 284
rect -603 281 -601 284
rect -570 281 -568 284
rect -546 282 -544 285
rect -522 282 -520 285
rect -496 282 -494 285
rect -420 282 -418 285
rect -394 282 -392 285
rect -370 282 -368 285
rect -653 269 -651 272
rect -629 269 -627 272
rect -603 270 -601 273
rect -346 281 -344 284
rect -311 281 -309 284
rect -257 281 -255 284
rect -233 282 -231 285
rect -209 282 -207 285
rect -183 282 -181 285
rect -677 261 -675 264
rect -653 261 -651 264
rect -629 261 -627 264
rect -807 248 -805 251
rect -781 246 -779 249
rect -757 247 -755 250
rect -653 255 -651 258
rect -603 257 -601 260
rect -570 257 -568 271
rect -546 269 -544 272
rect -522 269 -520 272
rect -496 269 -494 272
rect -420 269 -418 272
rect -394 269 -392 272
rect -370 269 -368 272
rect -546 257 -544 260
rect -522 257 -520 260
rect -496 258 -494 261
rect -420 258 -418 261
rect -629 254 -627 257
rect -653 247 -651 250
rect -807 240 -805 243
rect -708 244 -706 247
rect -629 246 -627 249
rect -603 248 -601 251
rect -570 249 -568 252
rect -546 249 -544 252
rect -522 249 -520 252
rect -394 257 -392 260
rect -370 257 -368 260
rect -346 257 -344 271
rect -151 281 -149 284
rect -127 282 -125 285
rect -103 282 -101 285
rect -77 282 -75 285
rect -394 249 -392 252
rect -370 249 -368 252
rect -346 249 -344 252
rect -546 243 -544 246
rect -496 245 -494 248
rect -420 245 -418 248
rect -311 246 -309 261
rect -257 257 -255 271
rect -233 269 -231 272
rect -209 269 -207 272
rect -183 269 -181 272
rect -233 257 -231 260
rect -209 257 -207 260
rect -183 258 -181 261
rect -257 249 -255 252
rect -233 249 -231 252
rect -209 249 -207 252
rect -151 257 -149 271
rect -127 269 -125 272
rect -103 269 -101 272
rect -77 269 -75 272
rect -127 257 -125 260
rect -103 257 -101 260
rect -77 258 -75 261
rect -151 249 -149 252
rect -127 249 -125 252
rect -103 249 -101 252
rect -603 240 -601 243
rect -522 242 -520 245
rect -394 242 -392 245
rect -370 243 -368 246
rect -546 235 -544 238
rect -522 234 -520 237
rect -496 236 -494 239
rect -420 236 -418 239
rect -394 234 -392 237
rect -370 235 -368 238
rect -233 243 -231 246
rect -183 245 -181 248
rect -209 242 -207 245
rect -127 243 -125 246
rect -77 245 -75 248
rect -496 228 -494 231
rect -420 228 -418 231
rect -311 233 -309 236
rect -233 235 -231 238
rect -209 234 -207 237
rect -183 236 -181 239
rect -103 242 -101 245
rect -127 235 -125 238
rect -103 234 -101 237
rect -77 236 -75 239
rect -183 228 -181 231
rect -77 228 -75 231
rect -56 208 -54 211
rect -32 209 -30 212
rect -8 209 -6 212
rect 18 209 20 212
rect -772 205 -769 207
rect -759 205 -744 207
rect -724 205 -721 207
rect -703 205 -700 207
rect -690 205 -672 207
rect -652 205 -649 207
rect -595 193 -592 195
rect -582 193 -567 195
rect -547 193 -544 195
rect -526 193 -523 195
rect -513 193 -495 195
rect -475 193 -472 195
rect -411 193 -408 195
rect -398 193 -383 195
rect -363 193 -360 195
rect -342 193 -339 195
rect -329 193 -311 195
rect -291 193 -288 195
rect -229 193 -226 195
rect -216 193 -201 195
rect -181 193 -178 195
rect -160 193 -157 195
rect -147 193 -129 195
rect -109 193 -106 195
rect -56 184 -54 198
rect -32 196 -30 199
rect -8 196 -6 199
rect 18 196 20 199
rect -32 184 -30 187
rect -8 184 -6 187
rect 18 185 20 188
rect -765 175 -762 177
rect -752 175 -737 177
rect -717 175 -714 177
rect -696 175 -693 177
rect -683 175 -665 177
rect -645 175 -642 177
rect -56 176 -54 179
rect -32 176 -30 179
rect -8 176 -6 179
rect -32 170 -30 173
rect 18 172 20 175
rect -8 169 -6 172
rect -588 163 -585 165
rect -575 163 -560 165
rect -540 163 -537 165
rect -519 163 -516 165
rect -506 163 -488 165
rect -468 163 -465 165
rect -404 163 -401 165
rect -391 163 -376 165
rect -356 163 -353 165
rect -335 163 -332 165
rect -322 163 -304 165
rect -284 163 -281 165
rect -222 163 -219 165
rect -209 163 -194 165
rect -174 163 -171 165
rect -153 163 -150 165
rect -140 163 -122 165
rect -102 163 -99 165
rect -732 151 -730 163
rect -660 151 -658 163
rect -32 162 -30 165
rect -8 161 -6 164
rect 18 163 20 166
rect 18 155 20 158
rect -758 141 -756 148
rect -689 141 -687 148
rect -555 139 -553 151
rect -483 139 -481 151
rect -371 139 -369 151
rect -299 139 -297 151
rect -189 139 -187 151
rect -117 139 -115 151
rect -758 128 -756 131
rect -732 128 -730 131
rect -689 128 -687 131
rect -660 128 -658 131
rect -581 129 -579 136
rect -512 129 -510 136
rect -397 129 -395 136
rect -328 129 -326 136
rect -215 129 -213 136
rect -146 129 -144 136
rect -66 130 -64 133
rect -42 131 -40 134
rect -18 131 -16 134
rect 8 131 10 134
rect -581 116 -579 119
rect -555 116 -553 119
rect -512 116 -510 119
rect -483 116 -481 119
rect -397 116 -395 119
rect -371 116 -369 119
rect -328 116 -326 119
rect -299 116 -297 119
rect -215 116 -213 119
rect -189 116 -187 119
rect -146 116 -144 119
rect -117 116 -115 119
rect -665 109 -663 112
rect -635 109 -633 112
rect -764 87 -762 91
rect -743 87 -741 91
rect -722 87 -720 91
rect -701 87 -699 91
rect -66 106 -64 120
rect -42 118 -40 121
rect -18 118 -16 121
rect 8 118 10 121
rect -42 106 -40 109
rect -18 106 -16 109
rect 8 107 10 110
rect -488 97 -486 100
rect -458 97 -456 100
rect -304 97 -302 100
rect -274 97 -272 100
rect -122 97 -120 100
rect -92 97 -90 100
rect -66 98 -64 101
rect -42 98 -40 101
rect -18 98 -16 101
rect -789 56 -787 59
rect -665 75 -663 89
rect -635 75 -633 89
rect -42 92 -40 95
rect 8 94 10 97
rect -18 91 -16 94
rect -42 84 -40 87
rect -18 83 -16 86
rect 8 85 10 88
rect 8 77 10 80
rect -488 63 -486 77
rect -458 63 -456 77
rect -304 63 -302 77
rect -274 63 -272 77
rect -122 63 -120 77
rect -92 63 -90 77
rect 66 63 68 66
rect -665 51 -663 55
rect -635 51 -633 55
rect -789 32 -787 46
rect -764 32 -762 47
rect -743 32 -741 47
rect -722 32 -720 47
rect -701 32 -699 47
rect -43 53 -41 56
rect -17 53 -15 56
rect 7 53 9 56
rect 31 52 33 55
rect -488 39 -486 43
rect -458 39 -456 43
rect -304 39 -302 43
rect -274 39 -272 43
rect -122 39 -120 43
rect -92 39 -90 43
rect -43 40 -41 43
rect -17 40 -15 43
rect 7 40 9 43
rect -419 35 -417 38
rect -398 35 -396 38
rect -377 35 -375 38
rect -641 27 -639 30
rect -620 27 -618 30
rect -599 27 -597 30
rect -578 27 -576 30
rect -789 9 -787 12
rect -764 9 -762 12
rect -743 9 -741 12
rect -722 9 -720 12
rect -701 9 -699 12
rect -43 29 -41 32
rect -492 12 -489 14
rect -479 12 -464 14
rect -444 12 -441 14
rect -694 -10 -692 -7
rect -674 -10 -672 -7
rect -641 -8 -639 7
rect -620 -8 -618 7
rect -599 -8 -597 7
rect -578 -8 -576 7
rect -419 0 -417 15
rect -398 0 -396 15
rect -377 0 -375 15
rect -240 18 -236 20
rect -216 18 -202 20
rect -182 18 -179 20
rect -17 28 -15 31
rect 7 28 9 31
rect 31 28 33 42
rect 66 28 68 43
rect -17 20 -15 23
rect 7 20 9 23
rect 31 20 33 23
rect -308 12 -305 14
rect -295 12 -280 14
rect -260 12 -257 14
rect -43 16 -41 19
rect -126 12 -123 14
rect -113 12 -98 14
rect -78 12 -75 14
rect -17 13 -15 16
rect 7 14 9 17
rect 66 15 68 18
rect -43 7 -41 10
rect -17 5 -15 8
rect 7 6 9 9
rect -856 -17 -854 -14
rect -822 -18 -820 -15
rect -801 -18 -799 -15
rect -780 -18 -778 -15
rect -759 -18 -757 -15
rect -856 -52 -854 -37
rect -822 -53 -820 -38
rect -801 -53 -799 -38
rect -780 -53 -778 -38
rect -759 -53 -757 -38
rect -694 -44 -692 -30
rect -674 -44 -672 -30
rect -856 -65 -854 -62
rect -476 -14 -474 -11
rect -456 -14 -454 -11
rect -240 -2 -236 0
rect -216 -2 -202 0
rect -182 -2 -179 0
rect -43 -1 -41 2
rect -292 -14 -290 -11
rect -272 -14 -270 -11
rect -110 -14 -108 -11
rect -90 -14 -88 -11
rect -419 -34 -417 -30
rect -398 -34 -396 -30
rect -377 -34 -375 -30
rect -476 -48 -474 -34
rect -456 -48 -454 -34
rect -292 -48 -290 -34
rect -272 -48 -270 -34
rect -110 -48 -108 -34
rect -90 -48 -88 -34
rect -53 -35 -51 -32
rect -29 -34 -27 -31
rect -5 -34 -3 -31
rect 21 -34 23 -31
rect -641 -52 -639 -48
rect -620 -52 -618 -48
rect -599 -52 -597 -48
rect -578 -52 -576 -48
rect -553 -59 -551 -56
rect -532 -59 -530 -56
rect -511 -59 -509 -56
rect -694 -68 -692 -64
rect -674 -68 -672 -64
rect -369 -56 -367 -53
rect -348 -56 -346 -53
rect -327 -56 -325 -53
rect -476 -72 -474 -68
rect -456 -71 -454 -68
rect -53 -59 -51 -45
rect -29 -47 -27 -44
rect -5 -47 -3 -44
rect 21 -47 23 -44
rect -29 -59 -27 -56
rect -5 -59 -3 -56
rect 21 -58 23 -55
rect -53 -67 -51 -64
rect -29 -67 -27 -64
rect -5 -67 -3 -64
rect -292 -72 -290 -68
rect -272 -72 -270 -68
rect -110 -72 -108 -68
rect -90 -72 -88 -68
rect -29 -73 -27 -70
rect 21 -71 23 -68
rect -638 -84 -636 -81
rect -617 -84 -615 -81
rect -596 -84 -594 -81
rect -822 -97 -820 -93
rect -801 -97 -799 -93
rect -780 -97 -778 -93
rect -759 -97 -757 -93
rect -731 -95 -729 -92
rect -710 -95 -708 -92
rect -689 -95 -687 -92
rect -668 -95 -666 -92
rect -812 -113 -809 -111
rect -789 -113 -775 -111
rect -755 -113 -751 -111
rect -553 -94 -551 -79
rect -532 -94 -530 -79
rect -511 -94 -509 -79
rect -369 -91 -367 -76
rect -348 -91 -346 -76
rect -327 -91 -325 -76
rect -5 -74 -3 -71
rect -29 -81 -27 -78
rect -216 -87 -214 -84
rect -190 -87 -188 -84
rect -166 -87 -164 -84
rect -5 -82 -3 -79
rect 21 -80 23 -77
rect -731 -130 -729 -115
rect -710 -130 -708 -115
rect -689 -130 -687 -115
rect -668 -130 -666 -115
rect -638 -119 -636 -104
rect -617 -119 -615 -104
rect -596 -119 -594 -104
rect -812 -133 -809 -131
rect -789 -133 -775 -131
rect -755 -133 -751 -131
rect -835 -162 -833 -159
rect -809 -162 -807 -159
rect -785 -162 -783 -159
rect -761 -163 -759 -160
rect -835 -175 -833 -172
rect -809 -175 -807 -172
rect -785 -175 -783 -172
rect -462 -95 -460 -92
rect -441 -95 -439 -92
rect -420 -95 -418 -92
rect -399 -95 -397 -92
rect -553 -128 -551 -124
rect -532 -128 -530 -124
rect -511 -128 -509 -124
rect -462 -130 -460 -115
rect -441 -130 -439 -115
rect -420 -130 -418 -115
rect -399 -130 -397 -115
rect -142 -88 -140 -85
rect 21 -88 23 -85
rect -216 -100 -214 -97
rect -190 -100 -188 -97
rect -166 -100 -164 -97
rect -216 -111 -214 -108
rect -190 -112 -188 -109
rect -166 -112 -164 -109
rect -142 -112 -140 -98
rect 21 -107 23 -104
rect -29 -114 -27 -111
rect -5 -113 -3 -110
rect -190 -120 -188 -117
rect -166 -120 -164 -117
rect -142 -120 -140 -117
rect 21 -115 23 -112
rect -369 -125 -367 -121
rect -348 -125 -346 -121
rect -327 -125 -325 -121
rect -216 -124 -214 -121
rect -29 -122 -27 -119
rect -5 -121 -3 -118
rect -190 -127 -188 -124
rect -166 -126 -164 -123
rect 21 -124 23 -121
rect -638 -153 -636 -149
rect -617 -153 -615 -149
rect -596 -153 -594 -149
rect -216 -133 -214 -130
rect -53 -128 -51 -125
rect -29 -128 -27 -125
rect -5 -128 -3 -125
rect -190 -135 -188 -132
rect -166 -134 -164 -131
rect -216 -141 -214 -138
rect -53 -147 -51 -133
rect -29 -136 -27 -133
rect -5 -136 -3 -133
rect 21 -137 23 -134
rect -29 -148 -27 -145
rect -5 -148 -3 -145
rect 21 -148 23 -145
rect -53 -160 -51 -157
rect -29 -161 -27 -158
rect -5 -161 -3 -158
rect 21 -161 23 -158
rect -150 -167 -147 -165
rect -137 -167 -122 -165
rect -102 -167 -99 -165
rect -835 -186 -833 -183
rect -809 -187 -807 -184
rect -785 -187 -783 -184
rect -761 -187 -759 -173
rect -731 -174 -729 -170
rect -710 -174 -708 -170
rect -689 -174 -687 -170
rect -668 -174 -666 -170
rect -462 -174 -460 -170
rect -441 -174 -439 -170
rect -420 -174 -418 -170
rect -399 -174 -397 -170
rect -634 -177 -630 -175
rect -610 -177 -596 -175
rect -576 -177 -573 -175
rect -809 -195 -807 -192
rect -785 -195 -783 -192
rect -761 -195 -759 -192
rect -835 -199 -833 -196
rect -809 -202 -807 -199
rect -785 -201 -783 -198
rect -634 -199 -630 -197
rect -610 -199 -596 -197
rect -576 -199 -573 -197
rect -835 -208 -833 -205
rect -809 -210 -807 -207
rect -785 -209 -783 -206
rect -835 -216 -833 -213
rect -761 -221 -758 -219
rect -738 -221 -723 -219
rect -713 -221 -710 -219
<< polycontact >>
rect -808 297 -804 301
rect -782 297 -778 301
rect -758 297 -754 301
rect -654 297 -650 301
rect -630 297 -626 301
rect -604 297 -600 301
rect -808 273 -804 277
rect -782 272 -778 276
rect -758 272 -754 276
rect -737 272 -733 276
rect -547 285 -543 289
rect -523 285 -519 289
rect -497 285 -493 289
rect -421 285 -417 289
rect -395 285 -391 289
rect -371 285 -367 289
rect -234 285 -230 289
rect -210 285 -206 289
rect -184 285 -180 289
rect -128 285 -124 289
rect -104 285 -100 289
rect -78 285 -74 289
rect -712 260 -708 264
rect -675 272 -671 276
rect -654 272 -650 276
rect -630 272 -626 276
rect -604 273 -600 277
rect -568 260 -564 264
rect -547 260 -543 264
rect -523 260 -519 264
rect -497 261 -493 265
rect -421 261 -417 265
rect -395 260 -391 264
rect -371 260 -367 264
rect -350 260 -346 264
rect -782 242 -778 246
rect -758 243 -754 247
rect -654 243 -650 247
rect -315 249 -311 253
rect -630 242 -626 246
rect -255 260 -251 264
rect -234 260 -230 264
rect -210 260 -206 264
rect -184 261 -180 265
rect -149 260 -145 264
rect -128 260 -124 264
rect -104 260 -100 264
rect -78 261 -74 265
rect -808 236 -804 240
rect -604 236 -600 240
rect -547 231 -543 235
rect -523 230 -519 234
rect -395 230 -391 234
rect -371 231 -367 235
rect -234 231 -230 235
rect -210 230 -206 234
rect -128 231 -124 235
rect -104 230 -100 234
rect -497 224 -493 228
rect -421 224 -417 228
rect -184 224 -180 228
rect -78 224 -74 228
rect -33 212 -29 216
rect -9 212 -5 216
rect 17 212 21 216
rect -756 207 -752 211
rect -687 207 -683 211
rect -579 195 -575 199
rect -510 195 -506 199
rect -395 195 -391 199
rect -326 195 -322 199
rect -213 195 -209 199
rect -144 195 -140 199
rect -54 187 -50 191
rect -33 187 -29 191
rect -9 187 -5 191
rect 17 188 21 192
rect -749 177 -745 181
rect -677 177 -673 181
rect -572 165 -568 169
rect -500 165 -496 169
rect -388 165 -384 169
rect -316 165 -312 169
rect -206 165 -202 169
rect -134 165 -130 169
rect -730 159 -726 163
rect -658 159 -654 163
rect -33 158 -29 162
rect -9 157 -5 161
rect 17 151 21 155
rect -762 144 -758 148
rect -693 144 -689 148
rect -553 147 -549 151
rect -481 147 -477 151
rect -369 147 -365 151
rect -297 147 -293 151
rect -187 147 -183 151
rect -115 147 -111 151
rect -585 132 -581 136
rect -516 132 -512 136
rect -401 132 -397 136
rect -332 132 -328 136
rect -219 132 -215 136
rect -150 132 -146 136
rect -43 134 -39 138
rect -19 134 -15 138
rect 7 134 11 138
rect -64 109 -60 113
rect -43 109 -39 113
rect -19 109 -15 113
rect 7 110 11 114
rect -669 78 -665 82
rect -633 78 -629 82
rect -43 80 -39 84
rect -19 79 -15 83
rect -492 66 -488 70
rect -456 66 -452 70
rect -308 66 -304 70
rect -272 66 -268 70
rect -126 66 -122 70
rect 7 73 11 77
rect -90 66 -86 70
rect -787 39 -783 43
rect -762 39 -758 43
rect -741 39 -737 43
rect -720 39 -716 43
rect -44 56 -40 60
rect -18 56 -14 60
rect 6 56 10 60
rect -699 39 -695 43
rect -476 14 -472 18
rect -44 32 -40 36
rect -18 31 -14 35
rect 6 31 10 35
rect 27 31 31 35
rect -213 20 -209 24
rect -639 -4 -635 0
rect -618 -4 -614 0
rect -597 -4 -593 0
rect -417 4 -413 8
rect -396 4 -392 8
rect -292 14 -288 18
rect 62 31 66 35
rect -110 14 -106 18
rect -375 4 -371 8
rect -576 -4 -572 0
rect -854 -49 -850 -45
rect -820 -49 -816 -45
rect -799 -49 -795 -45
rect -778 -49 -774 -45
rect -698 -41 -694 -37
rect -672 -41 -668 -37
rect -757 -49 -753 -45
rect -18 1 -14 5
rect 6 2 10 6
rect -213 -6 -209 -2
rect -44 -5 -40 -1
rect -30 -31 -26 -27
rect -6 -31 -2 -27
rect 20 -31 24 -27
rect -480 -45 -476 -41
rect -454 -45 -450 -41
rect -296 -45 -292 -41
rect -270 -45 -266 -41
rect -114 -45 -110 -41
rect -88 -45 -84 -41
rect -51 -56 -47 -52
rect -30 -56 -26 -52
rect -6 -56 -2 -52
rect 20 -55 24 -51
rect -782 -111 -778 -107
rect -551 -90 -547 -86
rect -530 -90 -526 -86
rect -509 -90 -505 -86
rect -367 -87 -363 -83
rect -346 -87 -342 -83
rect -325 -87 -321 -83
rect -217 -84 -213 -80
rect -191 -84 -187 -80
rect -167 -84 -163 -80
rect -30 -85 -26 -81
rect -729 -126 -725 -122
rect -708 -126 -704 -122
rect -687 -126 -683 -122
rect -636 -115 -632 -111
rect -615 -115 -611 -111
rect -594 -115 -590 -111
rect -666 -126 -662 -122
rect -782 -137 -778 -133
rect -836 -159 -832 -155
rect -810 -159 -806 -155
rect -786 -159 -782 -155
rect -460 -126 -456 -122
rect -439 -126 -435 -122
rect -418 -126 -414 -122
rect -6 -86 -2 -82
rect 20 -92 24 -88
rect -217 -108 -213 -104
rect -191 -109 -187 -105
rect -167 -109 -163 -105
rect -146 -109 -142 -105
rect 20 -104 24 -100
rect -30 -111 -26 -107
rect -6 -110 -2 -106
rect -397 -126 -393 -122
rect -191 -139 -187 -135
rect -167 -138 -163 -134
rect -217 -145 -213 -141
rect -51 -140 -47 -136
rect -30 -140 -26 -136
rect -6 -140 -2 -136
rect 20 -141 24 -137
rect -134 -165 -130 -161
rect -30 -165 -26 -161
rect -6 -165 -2 -161
rect 20 -165 24 -161
rect -836 -183 -832 -179
rect -810 -184 -806 -180
rect -786 -184 -782 -180
rect -765 -184 -761 -180
rect -607 -175 -603 -171
rect -607 -203 -603 -199
rect -810 -214 -806 -210
rect -786 -213 -782 -209
rect -836 -220 -832 -216
rect -730 -219 -726 -215
<< metal1 >>
rect -801 304 -790 307
rect -820 297 -808 300
rect -820 240 -817 297
rect -801 294 -798 304
rect -785 304 -623 307
rect -814 284 -812 287
rect -800 291 -798 294
rect -795 297 -782 300
rect -771 297 -758 300
rect -814 270 -811 284
rect -795 281 -792 297
rect -771 287 -768 297
rect -751 294 -748 304
rect -774 284 -768 287
rect -764 284 -762 287
rect -750 291 -748 294
rect -738 293 -734 304
rect -710 300 -706 304
rect -719 296 -695 300
rect -798 280 -792 281
rect -807 277 -801 279
rect -804 276 -801 277
rect -796 278 -792 280
rect -796 276 -795 278
rect -792 272 -782 275
rect -814 267 -812 270
rect -792 267 -789 272
rect -775 269 -772 284
rect -764 281 -761 284
rect -753 276 -748 277
rect -800 264 -789 267
rect -774 267 -772 269
rect -764 269 -761 276
rect -754 272 -748 276
rect -730 276 -726 283
rect -713 292 -709 296
rect -674 293 -670 304
rect -730 272 -720 276
rect -660 294 -657 304
rect -618 304 -581 307
rect -650 297 -637 300
rect -626 297 -613 300
rect -660 291 -658 294
rect -640 287 -637 297
rect -646 284 -644 287
rect -640 284 -634 287
rect -682 276 -678 283
rect -647 281 -644 284
rect -687 275 -678 276
rect -690 272 -678 275
rect -730 269 -726 272
rect -803 248 -800 260
rect -786 254 -783 264
rect -774 263 -771 267
rect -764 266 -762 269
rect -750 264 -749 267
rect -774 260 -766 263
rect -774 249 -772 252
rect -820 237 -808 240
rect -820 233 -817 237
rect -775 239 -772 249
rect -769 247 -766 260
rect -752 255 -749 264
rect -723 264 -720 272
rect -705 264 -701 272
rect -692 267 -687 272
rect -682 269 -678 272
rect -647 269 -644 276
rect -738 263 -734 264
rect -750 252 -749 255
rect -746 260 -734 263
rect -723 260 -712 264
rect -705 260 -695 264
rect -674 263 -670 264
rect -659 264 -658 267
rect -646 266 -644 269
rect -636 269 -633 284
rect -616 281 -613 297
rect -610 294 -607 304
rect -600 297 -588 300
rect -610 291 -608 294
rect -596 284 -594 287
rect -616 280 -610 281
rect -616 278 -612 280
rect -613 276 -612 278
rect -607 277 -601 279
rect -607 276 -604 277
rect -626 272 -616 275
rect -636 267 -634 269
rect -674 260 -662 263
rect -769 244 -758 247
rect -746 243 -743 260
rect -705 257 -701 260
rect -713 243 -709 247
rect -746 239 -695 243
rect -746 237 -743 239
rect -770 234 -743 237
rect -665 237 -662 260
rect -659 255 -656 264
rect -637 263 -634 267
rect -619 267 -616 272
rect -597 270 -594 284
rect -619 264 -608 267
rect -642 260 -634 263
rect -659 252 -658 255
rect -642 247 -639 260
rect -625 254 -622 264
rect -650 244 -639 247
rect -636 249 -634 252
rect -596 267 -594 270
rect -636 239 -633 249
rect -608 248 -605 260
rect -626 242 -620 246
rect -625 241 -620 242
rect -591 240 -588 297
rect -584 295 -581 304
rect -584 292 -516 295
rect -567 281 -563 292
rect -553 282 -550 292
rect -511 292 -403 295
rect -543 285 -530 288
rect -519 285 -506 288
rect -553 279 -551 282
rect -533 275 -530 285
rect -539 272 -537 275
rect -533 272 -527 275
rect -575 264 -571 271
rect -540 269 -537 272
rect -582 260 -571 264
rect -582 256 -579 260
rect -575 257 -571 260
rect -540 257 -537 264
rect -583 251 -578 256
rect -567 251 -563 252
rect -552 252 -551 255
rect -539 254 -537 257
rect -529 257 -526 272
rect -509 269 -506 285
rect -503 282 -500 292
rect -493 285 -481 288
rect -503 279 -501 282
rect -489 272 -487 275
rect -509 268 -503 269
rect -509 266 -505 268
rect -506 264 -505 266
rect -500 265 -494 267
rect -500 264 -497 265
rect -519 260 -509 263
rect -529 255 -527 257
rect -567 248 -555 251
rect -665 234 -638 237
rect -600 237 -588 240
rect -820 230 -798 233
rect -801 190 -798 230
rect -558 225 -555 248
rect -552 243 -549 252
rect -530 251 -527 255
rect -512 255 -509 260
rect -490 258 -487 272
rect -512 252 -501 255
rect -535 248 -527 251
rect -552 240 -551 243
rect -535 235 -532 248
rect -518 242 -515 252
rect -543 232 -532 235
rect -529 237 -527 240
rect -489 255 -487 258
rect -529 227 -526 237
rect -501 236 -498 248
rect -519 230 -513 234
rect -518 229 -513 230
rect -484 228 -481 285
rect -433 285 -421 288
rect -443 268 -438 269
rect -433 268 -430 285
rect -414 282 -411 292
rect -398 292 -203 295
rect -443 265 -430 268
rect -443 264 -438 265
rect -756 221 -708 225
rect -773 208 -769 212
rect -756 211 -752 221
rect -720 212 -716 218
rect -724 208 -716 212
rect -759 200 -744 204
rect -756 197 -752 200
rect -770 194 -752 197
rect -720 198 -716 208
rect -801 187 -788 190
rect -770 182 -766 194
rect -770 178 -762 182
rect -749 181 -745 185
rect -712 182 -708 221
rect -687 221 -636 225
rect -558 222 -531 225
rect -493 225 -481 228
rect -433 228 -430 265
rect -427 272 -425 275
rect -413 279 -411 282
rect -408 285 -395 288
rect -384 285 -371 288
rect -427 258 -424 272
rect -408 269 -405 285
rect -384 275 -381 285
rect -364 282 -361 292
rect -387 272 -381 275
rect -377 272 -375 275
rect -363 279 -361 282
rect -351 281 -347 292
rect -312 289 -308 292
rect -322 285 -298 289
rect -316 281 -312 285
rect -254 281 -250 292
rect -411 268 -405 269
rect -420 265 -414 267
rect -417 264 -414 265
rect -409 266 -405 268
rect -409 264 -408 266
rect -405 260 -395 263
rect -427 255 -425 258
rect -405 255 -402 260
rect -388 257 -385 272
rect -377 269 -374 272
rect -413 252 -402 255
rect -387 255 -385 257
rect -377 257 -374 264
rect -343 264 -339 271
rect -343 260 -327 264
rect -240 282 -237 292
rect -198 292 -97 295
rect -230 285 -217 288
rect -206 285 -193 288
rect -240 279 -238 282
rect -220 275 -217 285
rect -226 272 -224 275
rect -220 272 -214 275
rect -262 264 -258 271
rect -227 269 -224 272
rect -343 257 -339 260
rect -416 236 -413 248
rect -399 242 -396 252
rect -387 251 -384 255
rect -377 254 -375 257
rect -363 252 -362 255
rect -387 248 -379 251
rect -387 237 -385 240
rect -401 230 -395 234
rect -401 229 -396 230
rect -433 225 -421 228
rect -388 227 -385 237
rect -382 235 -379 248
rect -365 243 -362 252
rect -331 253 -327 260
rect -308 253 -304 261
rect -272 260 -258 264
rect -272 259 -267 260
rect -262 257 -258 260
rect -227 257 -224 264
rect -351 251 -347 252
rect -363 240 -362 243
rect -359 248 -347 251
rect -331 249 -315 253
rect -308 249 -298 253
rect -254 251 -250 252
rect -239 252 -238 255
rect -226 254 -224 257
rect -216 257 -213 272
rect -196 269 -193 285
rect -190 282 -187 292
rect -180 285 -168 288
rect -190 279 -188 282
rect -176 272 -174 275
rect -196 268 -190 269
rect -196 266 -192 268
rect -193 264 -192 266
rect -187 265 -181 267
rect -187 264 -184 265
rect -206 260 -196 263
rect -216 255 -214 257
rect -382 232 -371 235
rect -359 231 -356 248
rect -308 246 -304 249
rect -254 248 -242 251
rect -316 232 -312 236
rect -322 231 -298 232
rect -359 228 -298 231
rect -359 225 -356 228
rect -383 222 -356 225
rect -245 225 -242 248
rect -239 243 -236 252
rect -217 251 -214 255
rect -199 255 -196 260
rect -177 258 -174 272
rect -199 252 -188 255
rect -222 248 -214 251
rect -239 240 -238 243
rect -222 235 -219 248
rect -205 242 -202 252
rect -230 232 -219 235
rect -216 237 -214 240
rect -176 255 -174 258
rect -216 227 -213 237
rect -188 236 -185 248
rect -206 230 -200 234
rect -205 229 -200 230
rect -171 228 -168 285
rect -148 281 -144 292
rect -134 282 -131 292
rect -92 292 -49 295
rect -124 285 -111 288
rect -100 285 -87 288
rect -134 279 -132 282
rect -114 275 -111 285
rect -120 272 -118 275
rect -114 272 -108 275
rect -156 264 -152 271
rect -121 269 -118 272
rect -165 260 -152 264
rect -165 259 -160 260
rect -156 257 -152 260
rect -121 257 -118 264
rect -148 251 -144 252
rect -133 252 -132 255
rect -120 254 -118 257
rect -110 257 -107 272
rect -90 269 -87 285
rect -84 282 -81 292
rect -74 285 -62 288
rect -84 279 -82 282
rect -70 272 -68 275
rect -90 268 -84 269
rect -90 266 -86 268
rect -87 264 -86 266
rect -81 265 -75 267
rect -81 264 -78 265
rect -100 260 -90 263
rect -110 255 -108 257
rect -148 248 -136 251
rect -245 222 -218 225
rect -180 225 -168 228
rect -139 225 -136 248
rect -133 243 -130 252
rect -111 251 -108 255
rect -93 255 -90 260
rect -71 258 -68 272
rect -93 252 -82 255
rect -116 248 -108 251
rect -133 240 -132 243
rect -116 235 -113 248
rect -99 242 -96 252
rect -124 232 -113 235
rect -110 237 -108 240
rect -70 255 -68 258
rect -110 227 -107 237
rect -82 236 -79 248
rect -100 230 -94 234
rect -99 229 -94 230
rect -65 228 -62 285
rect -139 222 -112 225
rect -74 225 -62 228
rect -52 222 -49 292
rect -687 211 -683 221
rect -648 212 -644 218
rect -652 208 -644 212
rect -690 200 -672 204
rect -687 197 -683 200
rect -770 148 -766 178
rect -717 178 -708 182
rect -752 170 -737 174
rect -749 163 -745 170
rect -712 163 -708 178
rect -754 160 -733 163
rect -754 158 -751 160
rect -770 144 -762 148
rect -755 141 -751 158
rect -737 151 -733 160
rect -726 159 -713 163
rect -763 127 -759 131
rect -729 127 -725 131
rect -763 123 -750 127
rect -745 123 -719 127
rect -713 119 -708 158
rect -701 194 -683 197
rect -648 198 -644 208
rect -640 207 -636 221
rect -53 219 -2 222
rect -579 209 -531 213
rect -701 182 -697 194
rect -652 193 -648 196
rect -701 178 -693 182
rect -677 181 -673 185
rect -640 182 -636 202
rect -596 196 -592 200
rect -579 199 -575 209
rect -543 200 -539 206
rect -547 196 -539 200
rect -582 188 -567 192
rect -579 185 -575 188
rect -701 148 -697 178
rect -645 178 -636 182
rect -683 170 -665 174
rect -677 163 -673 170
rect -640 163 -636 178
rect -682 160 -661 163
rect -701 144 -693 148
rect -686 141 -682 158
rect -665 151 -661 160
rect -654 159 -636 163
rect -593 182 -575 185
rect -543 186 -539 196
rect -593 170 -589 182
rect -593 166 -585 170
rect -572 169 -568 173
rect -535 170 -531 209
rect -510 209 -459 213
rect -510 199 -506 209
rect -471 200 -467 206
rect -475 196 -467 200
rect -513 188 -495 192
rect -510 185 -506 188
rect -593 136 -589 166
rect -540 166 -531 170
rect -575 158 -560 162
rect -572 151 -568 158
rect -535 151 -531 166
rect -577 148 -556 151
rect -577 146 -574 148
rect -593 132 -585 136
rect -694 127 -690 131
rect -657 127 -653 131
rect -578 129 -574 146
rect -694 123 -678 127
rect -673 123 -647 127
rect -560 139 -556 148
rect -549 147 -536 151
rect -713 116 -685 119
rect -780 65 -777 92
rect -761 88 -744 91
rect -761 87 -757 88
rect -786 61 -777 65
rect -786 56 -783 61
rect -748 87 -744 88
rect -740 88 -723 91
rect -740 87 -736 88
rect -727 87 -723 88
rect -719 88 -702 91
rect -719 87 -715 88
rect -706 87 -702 88
rect -698 87 -694 92
rect -794 43 -790 46
rect -797 40 -790 43
rect -794 32 -790 40
rect -783 39 -779 43
rect -769 43 -765 47
rect -688 44 -685 116
rect -676 113 -652 117
rect -646 113 -622 117
rect -586 115 -582 119
rect -552 115 -548 119
rect -670 109 -666 113
rect -632 109 -628 113
rect -586 111 -573 115
rect -662 82 -658 89
rect -568 111 -542 115
rect -640 82 -636 89
rect -673 78 -669 82
rect -662 78 -653 82
rect -648 78 -636 82
rect -629 78 -625 82
rect -640 75 -636 78
rect -670 50 -666 55
rect -669 46 -666 50
rect -573 61 -568 110
rect -662 50 -658 55
rect -632 50 -628 55
rect -662 46 -628 50
rect -774 39 -765 43
rect -690 41 -685 44
rect -769 32 -765 39
rect -748 32 -744 39
rect -727 32 -723 39
rect -706 32 -702 39
rect -536 35 -531 146
rect -524 182 -506 185
rect -471 186 -467 196
rect -463 195 -459 209
rect -395 209 -347 213
rect -412 196 -408 200
rect -395 199 -391 209
rect -359 200 -355 206
rect -363 196 -355 200
rect -524 170 -520 182
rect -475 181 -471 184
rect -524 166 -516 170
rect -500 169 -496 173
rect -463 170 -459 190
rect -398 188 -383 192
rect -395 185 -391 188
rect -524 136 -520 166
rect -468 166 -459 170
rect -506 158 -488 162
rect -500 151 -496 158
rect -463 151 -459 166
rect -505 148 -484 151
rect -524 132 -516 136
rect -509 129 -505 146
rect -488 139 -484 148
rect -477 147 -459 151
rect -409 182 -391 185
rect -359 186 -355 196
rect -409 170 -405 182
rect -409 166 -401 170
rect -388 169 -384 173
rect -351 170 -347 209
rect -326 209 -275 213
rect -326 199 -322 209
rect -287 200 -283 206
rect -291 196 -283 200
rect -329 188 -311 192
rect -326 185 -322 188
rect -409 136 -405 166
rect -356 166 -347 170
rect -391 158 -376 162
rect -388 151 -384 158
rect -351 151 -347 166
rect -393 148 -372 151
rect -393 146 -390 148
rect -409 132 -401 136
rect -394 129 -390 146
rect -517 115 -513 119
rect -480 115 -476 119
rect -376 139 -372 148
rect -365 147 -352 151
rect -402 115 -398 119
rect -368 115 -364 119
rect -517 111 -501 115
rect -496 111 -470 115
rect -402 111 -389 115
rect -384 111 -358 115
rect -508 101 -475 105
rect -469 101 -445 105
rect -652 34 -565 35
rect -786 8 -782 12
rect -761 8 -757 12
rect -740 8 -736 12
rect -719 8 -715 12
rect -698 8 -694 12
rect -676 31 -550 34
rect -536 32 -511 35
rect -676 8 -673 31
rect -638 27 -634 31
rect -617 27 -613 31
rect -596 27 -592 31
rect -575 27 -571 31
rect -800 5 -673 8
rect -800 4 -688 5
rect -867 -10 -843 -9
rect -800 -10 -797 4
rect -676 -2 -673 5
rect -646 0 -642 7
rect -625 0 -621 7
rect -604 0 -600 7
rect -583 0 -579 7
rect -712 -5 -661 -2
rect -572 -4 -562 -1
rect -867 -13 -746 -10
rect -853 -17 -849 -13
rect -836 -14 -746 -13
rect -861 -45 -857 -37
rect -864 -49 -857 -45
rect -850 -49 -846 -45
rect -861 -52 -857 -49
rect -853 -63 -849 -62
rect -836 -100 -833 -14
rect -819 -18 -815 -14
rect -798 -18 -794 -14
rect -777 -18 -773 -14
rect -756 -18 -752 -14
rect -827 -45 -823 -38
rect -806 -45 -802 -38
rect -785 -45 -781 -38
rect -764 -45 -760 -38
rect -753 -49 -744 -46
rect -827 -53 -823 -50
rect -747 -53 -744 -49
rect -819 -94 -815 -93
rect -806 -94 -802 -93
rect -819 -97 -802 -94
rect -798 -94 -794 -93
rect -785 -94 -781 -93
rect -798 -97 -781 -94
rect -777 -94 -773 -93
rect -764 -94 -760 -93
rect -777 -97 -760 -94
rect -756 -94 -752 -93
rect -712 -76 -709 -5
rect -705 -6 -661 -5
rect -699 -10 -695 -6
rect -671 -10 -667 -6
rect -646 -8 -642 -5
rect -691 -36 -687 -30
rect -650 -14 -649 -11
rect -700 -41 -698 -37
rect -691 -40 -684 -36
rect -691 -44 -687 -40
rect -679 -40 -675 -30
rect -699 -69 -695 -64
rect -679 -69 -675 -64
rect -699 -73 -675 -69
rect -652 -55 -649 -14
rect -638 -49 -634 -48
rect -625 -49 -621 -48
rect -638 -52 -621 -49
rect -617 -49 -613 -48
rect -604 -49 -600 -48
rect -617 -52 -600 -49
rect -596 -49 -592 -48
rect -583 -49 -579 -48
rect -596 -52 -579 -49
rect -575 -49 -571 -48
rect -553 -51 -550 31
rect -514 -41 -511 32
rect -508 -5 -504 101
rect -493 97 -489 101
rect -455 97 -451 101
rect -485 70 -481 77
rect -463 70 -459 77
rect -496 66 -492 70
rect -485 66 -476 70
rect -471 66 -459 70
rect -452 66 -448 70
rect -493 40 -489 43
rect -492 35 -489 40
rect -485 37 -481 43
rect -476 45 -471 65
rect -463 63 -459 66
rect -389 61 -384 110
rect -455 37 -451 43
rect -430 39 -368 43
rect -497 20 -493 35
rect -485 34 -451 37
rect -416 35 -412 39
rect -395 35 -391 39
rect -374 35 -370 39
rect -493 15 -489 19
rect -476 18 -472 26
rect -440 19 -436 25
rect -444 15 -436 19
rect -479 7 -464 11
rect -476 2 -472 7
rect -503 -10 -448 -6
rect -440 -6 -436 15
rect -424 8 -420 15
rect -403 8 -399 15
rect -382 8 -378 15
rect -443 -10 -436 -6
rect -424 0 -420 3
rect -481 -14 -477 -10
rect -453 -14 -449 -10
rect -514 -43 -480 -41
rect -542 -45 -480 -43
rect -473 -44 -469 -34
rect -416 -31 -412 -30
rect -403 -31 -399 -30
rect -416 -34 -399 -31
rect -395 -31 -391 -30
rect -382 -31 -378 -30
rect -461 -41 -457 -34
rect -395 -35 -378 -31
rect -374 -31 -370 -30
rect -352 -38 -347 146
rect -340 182 -322 185
rect -287 186 -283 196
rect -279 195 -275 209
rect -213 209 -165 213
rect -230 196 -226 200
rect -213 199 -209 209
rect -177 200 -173 206
rect -181 196 -173 200
rect -340 170 -336 182
rect -291 181 -287 184
rect -340 166 -332 170
rect -316 169 -312 173
rect -279 170 -275 190
rect -216 188 -201 192
rect -213 185 -209 188
rect -340 136 -336 166
rect -284 166 -275 170
rect -322 158 -304 162
rect -316 151 -312 158
rect -279 151 -275 166
rect -321 148 -300 151
rect -340 132 -332 136
rect -325 129 -321 146
rect -304 139 -300 148
rect -293 147 -275 151
rect -227 182 -209 185
rect -177 186 -173 196
rect -227 170 -223 182
rect -227 166 -219 170
rect -206 169 -202 173
rect -169 170 -165 209
rect -144 209 -93 213
rect -144 199 -140 209
rect -105 200 -101 206
rect -109 196 -101 200
rect -147 188 -129 192
rect -144 185 -140 188
rect -227 136 -223 166
rect -174 166 -165 170
rect -209 158 -194 162
rect -206 151 -202 158
rect -169 151 -165 166
rect -211 148 -190 151
rect -211 146 -208 148
rect -227 132 -219 136
rect -212 129 -208 146
rect -333 115 -329 119
rect -296 115 -292 119
rect -194 139 -190 148
rect -183 147 -170 151
rect -158 182 -140 185
rect -105 186 -101 196
rect -97 195 -93 209
rect -53 208 -49 219
rect -39 209 -36 219
rect 3 219 14 222
rect -29 212 -16 215
rect -5 212 8 215
rect -39 206 -37 209
rect -19 202 -16 212
rect -25 199 -23 202
rect -19 199 -13 202
rect -61 191 -57 198
rect -26 196 -23 199
rect -158 170 -154 182
rect -109 181 -105 184
rect -135 173 -130 178
rect -158 166 -150 170
rect -134 169 -130 173
rect -97 170 -93 190
rect -71 187 -57 191
rect -39 187 -33 190
rect -71 186 -66 187
rect -61 184 -57 187
rect -26 184 -23 191
rect -53 178 -49 179
rect -38 179 -37 182
rect -25 181 -23 184
rect -15 184 -12 199
rect 5 196 8 212
rect 11 209 14 219
rect 21 212 33 215
rect 11 206 13 209
rect 25 199 27 202
rect 5 195 11 196
rect 5 193 9 195
rect 8 191 9 193
rect 14 192 20 194
rect 14 191 17 192
rect -5 187 5 190
rect -15 182 -13 184
rect -53 175 -41 178
rect -220 115 -216 119
rect -186 115 -182 119
rect -333 111 -317 115
rect -312 111 -286 115
rect -220 111 -207 115
rect -202 111 -176 115
rect -324 101 -291 105
rect -285 101 -261 105
rect -324 45 -320 101
rect -309 97 -305 101
rect -271 97 -267 101
rect -301 70 -297 77
rect -279 70 -275 77
rect -312 66 -308 70
rect -301 66 -292 70
rect -287 66 -275 70
rect -268 66 -264 70
rect -332 3 -329 31
rect -324 -6 -320 40
rect -309 38 -305 43
rect -308 34 -305 38
rect -301 37 -297 43
rect -292 45 -287 65
rect -279 63 -275 66
rect -207 61 -202 110
rect -271 37 -267 43
rect -301 34 -267 37
rect -313 20 -309 33
rect -309 15 -305 19
rect -292 18 -288 26
rect -256 19 -252 25
rect -213 24 -209 26
rect -178 25 -174 31
rect -182 21 -174 25
rect -260 15 -252 19
rect -295 7 -293 11
rect -288 7 -280 11
rect -256 -6 -252 15
rect -320 -10 -252 -6
rect -245 13 -236 17
rect -212 13 -202 17
rect -245 -3 -241 13
rect -212 6 -209 13
rect -216 1 -214 5
rect -209 1 -202 5
rect -245 -7 -236 -3
rect -178 -3 -174 21
rect -297 -14 -293 -10
rect -269 -14 -265 -10
rect -464 -44 -457 -41
rect -542 -46 -511 -45
rect -461 -48 -457 -44
rect -450 -45 -437 -41
rect -429 -43 -352 -40
rect -347 -40 -309 -39
rect -347 -41 -303 -40
rect -347 -43 -296 -41
rect -564 -55 -508 -51
rect -503 -55 -498 -51
rect -652 -58 -620 -55
rect -652 -62 -649 -58
rect -671 -73 -667 -64
rect -623 -69 -620 -58
rect -550 -59 -546 -55
rect -529 -59 -525 -55
rect -508 -59 -504 -55
rect -623 -72 -577 -69
rect -749 -94 -746 -76
rect -712 -79 -583 -76
rect -696 -87 -693 -79
rect -649 -80 -583 -79
rect -635 -84 -631 -80
rect -614 -84 -610 -80
rect -593 -84 -589 -80
rect -742 -91 -655 -87
rect -756 -97 -746 -94
rect -728 -95 -724 -91
rect -707 -95 -703 -91
rect -686 -95 -682 -91
rect -665 -95 -661 -91
rect -836 -103 -813 -100
rect -817 -106 -813 -103
rect -817 -110 -809 -106
rect -782 -107 -778 -105
rect -750 -106 -746 -97
rect -829 -127 -824 -122
rect -829 -143 -826 -127
rect -848 -146 -826 -143
rect -817 -134 -813 -110
rect -755 -110 -746 -106
rect -750 -111 -746 -110
rect -789 -118 -779 -114
rect -755 -118 -746 -114
rect -782 -121 -779 -118
rect -783 -126 -778 -121
rect -789 -130 -775 -126
rect -817 -138 -809 -134
rect -750 -134 -746 -118
rect -580 -102 -577 -72
rect -574 -87 -571 -63
rect -481 -73 -477 -68
rect -483 -77 -477 -73
rect -429 -49 -426 -43
rect -473 -71 -469 -68
rect -453 -71 -449 -68
rect -473 -74 -449 -71
rect -446 -52 -426 -49
rect -446 -77 -443 -52
rect -423 -71 -420 -43
rect -306 -44 -296 -43
rect -289 -44 -285 -34
rect -277 -41 -273 -34
rect -213 -41 -209 -6
rect -182 -7 -178 -3
rect -280 -44 -273 -41
rect -380 -51 -325 -48
rect -277 -48 -273 -44
rect -266 -45 -262 -41
rect -320 -51 -314 -48
rect -380 -52 -314 -51
rect -366 -56 -362 -52
rect -345 -56 -341 -52
rect -324 -56 -320 -52
rect -297 -73 -293 -68
rect -558 -86 -554 -79
rect -537 -86 -533 -79
rect -516 -86 -512 -79
rect -474 -80 -443 -77
rect -474 -81 -471 -80
rect -491 -84 -471 -81
rect -374 -83 -370 -76
rect -353 -83 -349 -76
rect -332 -83 -328 -76
rect -299 -77 -293 -73
rect -289 -73 -285 -68
rect -269 -73 -265 -68
rect -289 -77 -265 -73
rect -491 -86 -488 -84
rect -574 -90 -559 -87
rect -500 -90 -488 -86
rect -479 -90 -439 -87
rect -558 -94 -554 -91
rect -643 -111 -639 -104
rect -622 -111 -618 -104
rect -601 -111 -597 -104
rect -580 -105 -567 -102
rect -736 -122 -732 -115
rect -715 -122 -711 -115
rect -694 -122 -690 -115
rect -673 -122 -669 -115
rect -643 -119 -639 -116
rect -848 -156 -845 -146
rect -817 -148 -813 -138
rect -782 -141 -778 -137
rect -755 -138 -746 -134
rect -736 -130 -732 -127
rect -829 -152 -818 -149
rect -848 -159 -836 -156
rect -848 -216 -845 -159
rect -829 -162 -826 -152
rect -813 -152 -762 -149
rect -842 -172 -840 -169
rect -828 -165 -826 -162
rect -823 -159 -810 -156
rect -799 -159 -786 -156
rect -842 -186 -839 -172
rect -823 -175 -820 -159
rect -799 -169 -796 -159
rect -779 -162 -776 -152
rect -802 -172 -796 -169
rect -792 -172 -790 -169
rect -778 -165 -776 -162
rect -766 -163 -762 -152
rect -826 -176 -820 -175
rect -835 -179 -829 -177
rect -832 -180 -829 -179
rect -824 -178 -820 -176
rect -824 -180 -823 -178
rect -820 -184 -810 -181
rect -842 -189 -840 -186
rect -820 -189 -817 -184
rect -803 -187 -800 -172
rect -792 -175 -789 -172
rect -828 -192 -817 -189
rect -802 -189 -800 -187
rect -792 -187 -789 -180
rect -758 -180 -754 -173
rect -728 -171 -724 -170
rect -715 -171 -711 -170
rect -728 -174 -711 -171
rect -707 -171 -703 -170
rect -694 -171 -690 -170
rect -707 -174 -690 -171
rect -686 -171 -682 -170
rect -673 -171 -669 -170
rect -686 -174 -669 -171
rect -635 -150 -631 -149
rect -622 -150 -618 -149
rect -635 -153 -618 -150
rect -614 -150 -610 -149
rect -601 -150 -597 -149
rect -614 -153 -597 -150
rect -567 -123 -564 -105
rect -550 -125 -546 -124
rect -537 -125 -533 -124
rect -550 -128 -533 -125
rect -529 -125 -525 -124
rect -516 -125 -512 -124
rect -529 -128 -512 -125
rect -508 -125 -504 -124
rect -593 -154 -589 -149
rect -507 -154 -504 -130
rect -593 -156 -504 -154
rect -665 -171 -661 -170
rect -658 -157 -504 -156
rect -658 -159 -590 -157
rect -658 -171 -655 -159
rect -639 -168 -636 -159
rect -479 -160 -476 -90
rect -473 -91 -439 -90
rect -434 -91 -386 -87
rect -304 -84 -301 -78
rect -313 -87 -301 -84
rect -374 -91 -370 -88
rect -313 -91 -310 -87
rect -459 -95 -455 -91
rect -438 -95 -434 -91
rect -417 -95 -413 -91
rect -396 -95 -392 -91
rect -467 -122 -463 -115
rect -446 -122 -442 -115
rect -425 -122 -421 -115
rect -404 -122 -400 -115
rect -366 -122 -362 -121
rect -353 -122 -349 -121
rect -388 -127 -373 -124
rect -366 -125 -349 -122
rect -345 -122 -341 -121
rect -332 -122 -328 -121
rect -345 -125 -328 -122
rect -324 -122 -320 -121
rect -317 -94 -310 -91
rect -317 -122 -314 -94
rect -262 -97 -259 -46
rect -252 -105 -249 -53
rect -210 -77 -199 -74
rect -229 -84 -217 -81
rect -237 -100 -232 -99
rect -229 -100 -226 -84
rect -210 -87 -207 -77
rect -178 -74 -174 -8
rect -169 -42 -166 146
rect -158 136 -154 166
rect -102 166 -93 170
rect -140 158 -122 162
rect -134 151 -130 158
rect -97 151 -93 166
rect -139 148 -118 151
rect -158 132 -150 136
rect -143 129 -139 146
rect -122 139 -118 148
rect -111 147 -93 151
rect -44 152 -41 175
rect -38 170 -35 179
rect -16 178 -13 182
rect 2 182 5 187
rect 24 185 27 199
rect 2 179 13 182
rect -21 175 -13 178
rect -38 167 -37 170
rect -21 162 -18 175
rect -4 169 -1 179
rect -29 159 -18 162
rect -15 164 -13 167
rect 25 182 27 185
rect -15 154 -12 164
rect 13 163 16 175
rect 30 155 33 212
rect -44 149 -17 152
rect 21 152 33 155
rect -63 141 -12 144
rect -63 130 -59 141
rect -151 115 -147 119
rect -114 115 -110 119
rect -49 131 -46 141
rect -7 141 29 144
rect -39 134 -26 137
rect -15 134 -2 137
rect -49 128 -47 131
rect -29 124 -26 134
rect -35 121 -33 124
rect -29 121 -23 124
rect -151 111 -135 115
rect -130 111 -104 115
rect -71 113 -67 120
rect -36 118 -33 121
rect -77 109 -67 113
rect -49 109 -43 113
rect -71 106 -67 109
rect -36 106 -33 113
rect -142 101 -109 105
rect -103 101 -79 105
rect -142 -3 -138 101
rect -127 97 -123 101
rect -89 97 -85 101
rect -63 100 -59 101
rect -48 101 -47 104
rect -35 103 -33 106
rect -25 106 -22 121
rect -5 118 -2 134
rect 1 131 4 141
rect 11 134 23 137
rect 1 128 3 131
rect 15 121 17 124
rect -5 117 1 118
rect -5 115 -1 117
rect -2 113 -1 115
rect 4 114 10 116
rect 4 113 7 114
rect -15 109 -5 112
rect -25 104 -23 106
rect -63 97 -51 100
rect -119 70 -115 77
rect -54 78 -51 97
rect -48 92 -45 101
rect -26 100 -23 104
rect -8 104 -5 109
rect 14 107 17 121
rect -8 101 3 104
rect -31 97 -23 100
rect -48 89 -47 92
rect -31 84 -28 97
rect -14 91 -11 101
rect -39 81 -28 84
rect -25 86 -23 89
rect 15 104 17 107
rect -97 70 -93 77
rect -25 76 -22 86
rect 3 85 6 97
rect 20 77 23 134
rect -49 73 -27 74
rect -54 71 -27 73
rect 11 74 23 77
rect -130 66 -126 70
rect -119 66 -110 70
rect -105 66 -93 70
rect -86 66 -82 70
rect -127 40 -123 43
rect -126 35 -123 40
rect -110 49 -105 65
rect -97 63 -93 66
rect -37 63 -26 66
rect -119 37 -115 43
rect -89 37 -85 43
rect -131 20 -127 35
rect -119 34 -85 37
rect -56 56 -44 59
rect -56 32 -53 56
rect -37 53 -34 63
rect 26 66 29 141
rect 47 68 79 71
rect 47 66 50 68
rect 55 67 79 68
rect -21 63 50 66
rect -59 27 -53 32
rect -127 15 -123 19
rect -110 18 -106 26
rect -74 19 -70 25
rect -78 15 -70 19
rect -113 7 -98 11
rect -110 2 -106 7
rect -74 -6 -70 15
rect -56 -1 -53 27
rect -50 43 -48 46
rect -36 50 -34 53
rect -31 56 -18 59
rect -7 56 6 59
rect -50 29 -47 43
rect -31 40 -28 56
rect -7 46 -4 56
rect 13 53 16 63
rect -10 43 -4 46
rect 0 43 2 46
rect 14 50 16 53
rect 26 52 30 63
rect -34 39 -28 40
rect -43 36 -37 38
rect -40 35 -37 36
rect -32 37 -28 39
rect -32 35 -31 37
rect -28 31 -18 34
rect -50 26 -48 29
rect -28 26 -25 31
rect -11 28 -8 43
rect 0 40 3 43
rect 11 35 16 36
rect -36 23 -25 26
rect -10 26 -8 28
rect 0 28 3 35
rect 10 31 16 35
rect 34 35 38 42
rect 34 30 43 35
rect 34 28 38 30
rect -39 7 -36 19
rect -22 13 -19 23
rect -10 22 -7 26
rect 0 25 2 28
rect 14 23 15 26
rect -10 19 -2 22
rect -10 8 -8 11
rect -56 -4 -44 -1
rect -11 -2 -8 8
rect -5 6 -2 19
rect 12 14 15 23
rect 26 22 30 23
rect 14 11 15 14
rect 18 19 30 22
rect -5 3 6 6
rect -138 -8 -70 -6
rect 18 -4 21 19
rect -6 -7 21 -4
rect -142 -10 -70 -8
rect -115 -14 -111 -10
rect -87 -14 -83 -10
rect -169 -45 -114 -42
rect -107 -44 -103 -34
rect 47 -20 50 63
rect 61 63 65 67
rect 69 35 73 43
rect 53 31 62 35
rect 69 31 79 35
rect 53 30 58 31
rect 69 28 73 31
rect 61 14 65 18
rect 55 10 79 14
rect 55 9 60 10
rect -50 -24 1 -21
rect -95 -41 -91 -34
rect -50 -35 -46 -24
rect -98 -44 -91 -41
rect -169 -57 -166 -45
rect -95 -48 -91 -44
rect -84 -45 -71 -41
rect -36 -34 -33 -24
rect 12 -21 50 -20
rect 6 -23 50 -21
rect 6 -24 17 -23
rect 12 -25 17 -24
rect -26 -31 -13 -28
rect -2 -31 11 -28
rect -36 -37 -34 -34
rect -16 -41 -13 -31
rect -22 -44 -20 -41
rect -16 -44 -10 -41
rect -115 -73 -111 -68
rect -194 -77 -143 -74
rect -237 -103 -226 -100
rect -237 -104 -232 -103
rect -324 -125 -314 -122
rect -311 -108 -249 -105
rect -572 -163 -476 -160
rect -467 -130 -463 -127
rect -611 -167 -603 -164
rect -665 -174 -655 -171
rect -648 -170 -636 -168
rect -648 -171 -630 -170
rect -758 -185 -750 -180
rect -648 -182 -645 -171
rect -639 -174 -630 -171
rect -607 -171 -603 -167
rect -572 -170 -568 -163
rect -576 -174 -568 -170
rect -734 -185 -645 -182
rect -639 -182 -630 -178
rect -606 -181 -596 -178
rect -758 -187 -754 -185
rect -831 -208 -828 -196
rect -814 -202 -811 -192
rect -802 -193 -799 -189
rect -792 -190 -790 -187
rect -778 -192 -777 -189
rect -802 -196 -794 -193
rect -802 -207 -800 -204
rect -816 -214 -810 -210
rect -816 -215 -811 -214
rect -848 -219 -836 -216
rect -803 -217 -800 -207
rect -797 -209 -794 -196
rect -780 -201 -777 -192
rect -766 -193 -762 -192
rect -778 -204 -777 -201
rect -774 -196 -762 -193
rect -774 -201 -771 -196
rect -734 -201 -731 -185
rect -774 -204 -731 -201
rect -797 -212 -786 -209
rect -774 -219 -771 -204
rect -728 -208 -723 -206
rect -798 -222 -771 -219
rect -766 -214 -762 -208
rect -729 -211 -723 -208
rect -766 -218 -758 -214
rect -730 -215 -726 -211
rect -709 -214 -705 -185
rect -639 -200 -635 -182
rect -606 -184 -603 -181
rect -606 -192 -603 -189
rect -610 -196 -596 -192
rect -639 -204 -630 -200
rect -572 -200 -568 -174
rect -774 -226 -769 -225
rect -766 -226 -762 -218
rect -713 -218 -705 -214
rect -606 -213 -603 -203
rect -576 -204 -568 -200
rect -572 -210 -568 -204
rect -565 -169 -470 -166
rect -565 -213 -562 -169
rect -473 -179 -470 -169
rect -459 -171 -455 -170
rect -446 -171 -442 -170
rect -459 -174 -442 -171
rect -438 -171 -434 -170
rect -425 -171 -421 -170
rect -438 -174 -421 -171
rect -417 -171 -413 -170
rect -404 -171 -400 -170
rect -417 -174 -400 -171
rect -396 -171 -392 -170
rect -385 -179 -382 -127
rect -376 -128 -373 -127
rect -311 -128 -308 -108
rect -376 -131 -308 -128
rect -229 -141 -226 -103
rect -223 -97 -221 -94
rect -209 -90 -207 -87
rect -204 -84 -191 -81
rect -180 -84 -167 -81
rect -223 -111 -220 -97
rect -204 -100 -201 -84
rect -180 -94 -177 -84
rect -160 -87 -157 -77
rect -183 -97 -177 -94
rect -173 -97 -171 -94
rect -159 -90 -157 -87
rect -147 -88 -143 -77
rect -117 -77 -111 -73
rect -58 -52 -54 -45
rect -23 -47 -20 -44
rect -66 -56 -54 -52
rect -66 -60 -63 -56
rect -58 -59 -54 -56
rect -23 -59 -20 -52
rect -67 -65 -62 -60
rect -50 -65 -46 -64
rect -35 -64 -34 -61
rect -22 -62 -20 -59
rect -12 -59 -9 -44
rect 8 -47 11 -31
rect 14 -34 17 -25
rect 24 -31 36 -28
rect 14 -37 16 -34
rect 28 -44 30 -41
rect 8 -48 14 -47
rect 8 -50 12 -48
rect 11 -52 12 -50
rect 17 -51 23 -49
rect 17 -52 20 -51
rect -2 -56 8 -53
rect -12 -61 -10 -59
rect -50 -68 -38 -65
rect -107 -73 -103 -68
rect -87 -73 -83 -68
rect -107 -77 -83 -73
rect -114 -83 -111 -77
rect -41 -83 -38 -68
rect -35 -73 -32 -64
rect -13 -65 -10 -61
rect 5 -61 8 -56
rect 27 -58 30 -44
rect 5 -64 16 -61
rect -18 -68 -10 -65
rect -35 -76 -34 -73
rect -18 -81 -15 -68
rect -1 -74 2 -64
rect -114 -86 -38 -83
rect -26 -84 -15 -81
rect -12 -79 -10 -76
rect 28 -61 30 -58
rect -207 -101 -201 -100
rect -216 -104 -210 -102
rect -213 -105 -210 -104
rect -205 -103 -201 -101
rect -205 -105 -204 -103
rect -201 -109 -191 -106
rect -223 -114 -221 -111
rect -201 -114 -198 -109
rect -184 -112 -181 -97
rect -173 -100 -170 -97
rect -209 -117 -198 -114
rect -183 -114 -181 -112
rect -173 -112 -170 -105
rect -139 -105 -135 -98
rect -139 -109 -125 -105
rect -139 -112 -135 -109
rect -130 -110 -125 -109
rect -212 -133 -209 -121
rect -195 -127 -192 -117
rect -183 -118 -180 -114
rect -173 -115 -171 -112
rect -159 -117 -158 -114
rect -183 -121 -175 -118
rect -183 -132 -181 -129
rect -197 -139 -191 -135
rect -197 -140 -192 -139
rect -229 -144 -217 -141
rect -184 -142 -181 -132
rect -178 -134 -175 -121
rect -161 -126 -158 -117
rect -147 -118 -143 -117
rect -159 -129 -158 -126
rect -155 -121 -143 -118
rect -178 -137 -167 -134
rect -155 -142 -152 -121
rect -114 -142 -111 -86
rect -41 -91 -38 -86
rect -12 -89 -9 -79
rect 16 -80 19 -68
rect -2 -86 4 -82
rect -1 -87 4 -86
rect 33 -88 36 -31
rect -41 -94 -14 -91
rect 24 -91 36 -88
rect -41 -101 -14 -98
rect -41 -124 -38 -101
rect -26 -111 -15 -108
rect -66 -131 -61 -126
rect -50 -127 -38 -124
rect -35 -119 -34 -116
rect -50 -128 -46 -127
rect -65 -136 -62 -131
rect -35 -128 -32 -119
rect -18 -124 -15 -111
rect -12 -113 -9 -103
rect 24 -104 36 -101
rect -1 -106 4 -105
rect -2 -110 4 -106
rect -12 -116 -10 -113
rect -18 -127 -10 -124
rect -35 -131 -34 -128
rect -22 -133 -20 -130
rect -13 -131 -10 -127
rect -1 -128 2 -118
rect 16 -124 19 -112
rect -58 -136 -54 -133
rect -65 -140 -54 -136
rect -155 -144 -111 -142
rect -179 -145 -111 -144
rect -179 -147 -151 -145
rect -154 -160 -151 -147
rect -58 -147 -54 -140
rect -23 -140 -20 -133
rect -12 -133 -10 -131
rect 5 -131 16 -128
rect -135 -156 -130 -151
rect -154 -164 -147 -160
rect -134 -161 -130 -156
rect -98 -160 -94 -154
rect -23 -148 -20 -145
rect -12 -148 -9 -133
rect 5 -136 8 -131
rect 28 -134 30 -131
rect -2 -139 8 -136
rect 11 -142 12 -140
rect 8 -144 12 -142
rect 17 -141 20 -140
rect 17 -143 23 -141
rect 8 -145 14 -144
rect -154 -178 -151 -164
rect -102 -164 -94 -160
rect -98 -168 -94 -164
rect -50 -168 -46 -157
rect -36 -158 -34 -155
rect -22 -151 -20 -148
rect -16 -151 -10 -148
rect -36 -168 -33 -158
rect -16 -161 -13 -151
rect 8 -161 11 -145
rect 27 -148 30 -134
rect -26 -164 -13 -161
rect -2 -164 11 -161
rect 14 -158 16 -155
rect 28 -151 30 -148
rect -137 -172 -122 -168
rect -98 -171 1 -168
rect -134 -178 -130 -172
rect -98 -178 -94 -171
rect 14 -168 17 -158
rect 33 -161 36 -104
rect 24 -164 36 -161
rect 6 -171 17 -168
rect 12 -173 17 -171
rect -473 -182 -382 -179
rect -606 -216 -562 -213
rect -738 -226 -723 -222
rect -774 -229 -762 -226
rect -774 -230 -769 -229
rect -766 -232 -762 -229
rect -730 -232 -726 -226
rect -709 -232 -705 -218
<< m2contact >>
rect -82 109 -77 114
<< metal2 >>
rect -764 281 -739 284
rect -742 277 -739 281
rect -669 281 -644 284
rect -669 277 -666 281
rect -799 272 -796 275
rect -753 272 -748 277
rect -612 272 -609 275
rect -799 269 -749 272
rect -659 269 -609 272
rect -814 237 -811 248
rect -799 246 -796 269
rect -799 243 -787 246
rect -814 234 -775 237
rect -763 237 -760 255
rect -648 237 -645 255
rect -612 246 -609 269
rect -562 269 -537 272
rect -562 265 -559 269
rect -377 269 -352 272
rect -355 265 -352 269
rect -249 269 -224 272
rect -249 265 -246 269
rect -505 260 -502 263
rect -552 257 -502 260
rect -625 243 -609 246
rect -625 241 -620 243
rect -770 234 -638 237
rect -597 237 -594 248
rect -633 234 -554 237
rect -557 225 -554 234
rect -541 225 -538 243
rect -505 234 -502 257
rect -412 260 -409 263
rect -143 269 -118 272
rect -143 265 -140 269
rect -192 260 -189 263
rect -86 260 -83 263
rect -412 257 -362 260
rect -239 257 -189 260
rect -133 257 -83 260
rect -518 231 -502 234
rect -518 229 -513 231
rect -557 222 -531 225
rect -490 225 -487 236
rect -427 225 -424 236
rect -412 234 -409 257
rect -412 231 -396 234
rect -401 229 -396 231
rect -526 222 -388 225
rect -376 225 -373 243
rect -228 225 -225 243
rect -192 234 -189 257
rect -205 231 -189 234
rect -205 229 -200 231
rect -383 222 -218 225
rect -177 225 -174 236
rect -122 225 -119 243
rect -86 234 -83 257
rect -99 231 -83 234
rect -99 229 -94 231
rect -213 222 -112 225
rect -71 225 -68 236
rect -107 222 -68 225
rect -635 202 -620 207
rect -783 185 -754 190
rect -759 163 -754 185
rect -750 127 -745 185
rect -708 158 -687 163
rect -678 127 -673 185
rect -749 117 -746 122
rect -725 119 -682 122
rect -725 117 -722 119
rect -749 114 -722 117
rect -776 92 -698 97
rect -780 77 -777 92
rect -823 74 -777 77
rect -823 -3 -820 74
rect -806 52 -803 63
rect -809 49 -803 52
rect -809 36 -806 49
rect -777 48 -704 51
rect -777 44 -774 48
rect -749 44 -746 48
rect -728 44 -725 48
rect -707 44 -704 48
rect -809 33 -803 36
rect -853 -6 -820 -3
rect -868 -72 -864 -50
rect -853 -63 -850 -6
rect -806 -7 -803 33
rect -756 5 -753 39
rect -756 2 -739 5
rect -742 -4 -739 2
rect -735 3 -732 39
rect -714 3 -711 39
rect -735 0 -718 3
rect -714 0 -689 3
rect -721 -4 -718 0
rect -742 -7 -725 -4
rect -721 -7 -696 -4
rect -815 -10 -803 -7
rect -815 -45 -812 -10
rect -728 -11 -725 -7
rect -728 -14 -703 -11
rect -706 -22 -703 -14
rect -699 -15 -696 -7
rect -692 -8 -689 0
rect -685 -1 -682 119
rect -678 82 -673 122
rect -625 82 -620 202
rect -161 201 -158 222
rect -48 196 -23 199
rect -458 190 -443 195
rect -274 190 -259 195
rect -92 190 -77 195
rect -48 192 -45 196
rect -609 173 -577 178
rect -582 151 -577 173
rect -573 115 -568 173
rect -531 146 -510 151
rect -501 115 -496 173
rect -652 68 -649 77
rect -501 70 -496 110
rect -448 70 -443 190
rect -427 173 -393 178
rect -398 151 -393 173
rect -389 115 -384 173
rect -347 146 -326 151
rect -317 140 -312 173
rect -277 140 -272 141
rect -317 137 -272 140
rect -317 115 -312 137
rect -277 136 -272 137
rect -317 70 -312 110
rect -264 70 -259 190
rect -245 173 -211 178
rect -216 151 -211 173
rect -207 115 -202 173
rect -165 146 -144 151
rect -135 115 -130 178
rect -135 70 -130 110
rect -82 114 -77 190
rect -39 187 -34 192
rect 9 187 12 190
rect -38 184 12 187
rect -27 152 -24 170
rect 9 161 12 184
rect 0 158 12 161
rect -27 149 -17 152
rect 24 152 27 163
rect -12 149 27 152
rect -58 118 -33 121
rect -58 114 -55 118
rect -49 109 -44 114
rect -1 109 2 112
rect -82 70 -77 109
rect -49 106 2 109
rect -37 74 -34 92
rect -1 83 2 106
rect 14 90 17 149
rect -10 80 2 83
rect -37 71 -27 74
rect 14 74 17 85
rect -22 71 17 74
rect -568 56 -427 61
rect -384 56 -245 61
rect -202 56 -61 61
rect -476 31 -471 40
rect -523 26 -476 29
rect -647 4 -579 7
rect -647 0 -644 4
rect -624 0 -621 4
rect -603 0 -600 4
rect -582 0 -579 4
rect -523 0 -520 26
rect -430 8 -427 56
rect -412 31 -332 34
rect -292 31 -287 40
rect -412 8 -409 31
rect -295 27 -292 29
rect -370 24 -292 27
rect -402 12 -379 15
rect -402 8 -399 12
rect -382 8 -379 12
rect -370 8 -367 24
rect -342 8 -293 11
rect -430 5 -425 8
rect -685 -4 -647 -1
rect -557 -4 -520 0
rect -481 -3 -477 2
rect -424 -1 -420 3
rect -403 -1 -399 3
rect -424 -4 -399 -1
rect -692 -9 -652 -8
rect -692 -11 -655 -9
rect -634 -11 -631 -5
rect -634 -14 -627 -11
rect -699 -18 -660 -15
rect -706 -25 -667 -22
rect -663 -23 -660 -18
rect -670 -29 -667 -25
rect -794 -34 -717 -31
rect -670 -32 -647 -29
rect -794 -45 -791 -34
rect -785 -41 -761 -38
rect -785 -45 -782 -41
rect -764 -45 -761 -41
rect -720 -43 -717 -34
rect -663 -41 -659 -36
rect -841 -49 -828 -46
rect -827 -54 -824 -50
rect -806 -54 -803 -50
rect -785 -54 -782 -50
rect -827 -57 -782 -54
rect -868 -75 -811 -72
rect -814 -97 -811 -75
rect -814 -100 -780 -97
rect -773 -98 -770 -50
rect -705 -81 -702 -41
rect -650 -46 -647 -32
rect -652 -49 -647 -46
rect -652 -59 -649 -49
rect -630 -51 -627 -14
rect -630 -54 -618 -51
rect -652 -62 -625 -59
rect -628 -74 -625 -62
rect -621 -67 -618 -54
rect -613 -59 -610 -5
rect -592 -9 -589 -5
rect -592 -12 -521 -9
rect -524 -14 -521 -12
rect -524 -17 -465 -14
rect -519 -41 -512 -38
rect -468 -40 -465 -17
rect -613 -62 -575 -59
rect -621 -70 -571 -67
rect -628 -77 -578 -74
rect -773 -101 -742 -98
rect -745 -123 -742 -101
rect -720 -99 -717 -81
rect -705 -84 -585 -81
rect -720 -102 -700 -99
rect -736 -118 -712 -115
rect -736 -122 -733 -118
rect -715 -122 -712 -118
rect -703 -122 -700 -102
rect -694 -118 -670 -115
rect -694 -122 -691 -118
rect -673 -122 -670 -118
rect -660 -122 -657 -84
rect -643 -107 -598 -104
rect -643 -111 -640 -107
rect -622 -111 -619 -107
rect -601 -111 -598 -107
rect -588 -111 -585 -84
rect -581 -116 -578 -77
rect -574 -109 -571 -70
rect -547 -79 -544 -48
rect -515 -66 -512 -41
rect -427 -45 -394 -42
rect -427 -51 -424 -45
rect -445 -54 -424 -51
rect -515 -69 -502 -66
rect -566 -82 -544 -79
rect -566 -100 -563 -82
rect -547 -86 -544 -82
rect -536 -82 -514 -79
rect -536 -86 -533 -82
rect -517 -86 -514 -82
rect -505 -86 -502 -69
rect -445 -79 -442 -54
rect -397 -56 -394 -45
rect -404 -59 -394 -56
rect -473 -82 -442 -79
rect -493 -85 -470 -82
rect -557 -95 -554 -91
rect -538 -95 -535 -91
rect -557 -98 -535 -95
rect -524 -95 -521 -91
rect -493 -95 -490 -85
rect -524 -98 -490 -95
rect -423 -100 -420 -76
rect -397 -90 -394 -59
rect -390 -83 -387 3
rect -342 -6 -337 8
rect -248 9 -245 56
rect -110 31 -105 44
rect -208 26 -110 31
rect -248 6 -209 9
rect -327 -2 -280 1
rect -363 -43 -352 -40
rect -363 -83 -360 -43
rect -325 -46 -322 -11
rect -283 -40 -280 -2
rect -110 -27 -107 -3
rect -253 -30 -107 -27
rect -253 -41 -250 -30
rect -257 -44 -250 -41
rect -208 -44 -103 -41
rect -66 -45 -61 56
rect 0 40 25 43
rect 22 36 25 40
rect -35 31 -32 34
rect 11 31 16 36
rect 38 34 43 35
rect 53 34 58 35
rect 38 31 58 34
rect -35 28 15 31
rect 38 30 43 31
rect 53 30 58 31
rect -50 -4 -47 7
rect -35 5 -32 28
rect -35 2 -23 5
rect -50 -7 -11 -4
rect 1 -4 4 14
rect -6 -7 4 -4
rect -314 -53 -253 -50
rect -71 -50 -66 -46
rect -248 -53 -66 -50
rect -45 -47 -20 -44
rect -45 -51 -42 -47
rect -353 -79 -328 -76
rect -353 -83 -349 -79
rect -332 -83 -328 -79
rect -314 -83 -311 -53
rect 12 -56 15 -53
rect -264 -60 -170 -57
rect -264 -82 -261 -60
rect -390 -86 -375 -83
rect -397 -93 -379 -90
rect -562 -105 -452 -102
rect -574 -112 -486 -109
rect -745 -126 -737 -123
rect -777 -145 -743 -142
rect -792 -175 -767 -172
rect -770 -179 -767 -175
rect -746 -176 -743 -145
rect -723 -148 -720 -127
rect -715 -131 -712 -127
rect -694 -131 -691 -127
rect -715 -134 -691 -131
rect -681 -139 -678 -127
rect -630 -132 -627 -116
rect -611 -125 -608 -116
rect -581 -119 -550 -116
rect -611 -128 -569 -125
rect -630 -135 -579 -132
rect -681 -141 -583 -139
rect -567 -141 -564 -128
rect -553 -130 -550 -119
rect -489 -123 -486 -112
rect -455 -122 -452 -105
rect -434 -103 -420 -100
rect -382 -99 -379 -93
rect -374 -92 -370 -88
rect -354 -92 -349 -88
rect -374 -95 -349 -92
rect -316 -87 -311 -83
rect -307 -85 -261 -82
rect -342 -92 -337 -88
rect -307 -92 -304 -85
rect -342 -95 -304 -92
rect -382 -102 -264 -99
rect -434 -122 -431 -103
rect -255 -106 -252 -60
rect -35 -59 15 -56
rect -24 -91 -21 -73
rect 12 -82 15 -59
rect -1 -85 15 -82
rect -1 -87 4 -85
rect -24 -94 -14 -91
rect 27 -91 30 -80
rect -9 -94 30 -91
rect -173 -100 -148 -97
rect -13 -98 -10 -94
rect -151 -104 -148 -100
rect -24 -101 -14 -98
rect -310 -109 -252 -106
rect -208 -109 -205 -106
rect -426 -118 -400 -115
rect -426 -122 -423 -118
rect -403 -122 -400 -118
rect -489 -126 -468 -123
rect -553 -133 -514 -130
rect -517 -134 -514 -133
rect -467 -131 -464 -127
rect -446 -131 -443 -127
rect -425 -131 -422 -127
rect -467 -134 -422 -131
rect -413 -131 -410 -127
rect -310 -131 -307 -109
rect -208 -112 -158 -109
rect -130 -110 -125 -105
rect -413 -134 -307 -131
rect -517 -135 -500 -134
rect -517 -137 -472 -135
rect -503 -138 -472 -137
rect -413 -138 -410 -134
rect -475 -141 -410 -138
rect -681 -142 -564 -141
rect -586 -144 -564 -142
rect -223 -144 -220 -133
rect -208 -135 -205 -112
rect -208 -138 -192 -135
rect -197 -140 -192 -138
rect -223 -147 -184 -144
rect -172 -144 -169 -126
rect -179 -147 -169 -144
rect -723 -151 -540 -148
rect -130 -148 -127 -110
rect -24 -119 -21 -101
rect -9 -101 30 -98
rect -1 -107 4 -105
rect -1 -110 15 -107
rect 12 -133 15 -110
rect 27 -112 30 -101
rect -35 -136 15 -133
rect 12 -139 15 -136
rect -45 -145 -42 -141
rect -45 -148 -20 -145
rect -135 -151 -127 -148
rect -135 -156 -130 -151
rect -746 -179 -640 -176
rect -827 -184 -824 -181
rect -827 -187 -777 -184
rect -755 -185 -750 -180
rect -842 -219 -839 -208
rect -827 -210 -824 -187
rect -753 -188 -750 -185
rect -643 -185 -640 -179
rect -643 -188 -607 -185
rect -753 -191 -722 -188
rect -827 -213 -811 -210
rect -816 -215 -811 -213
rect -842 -222 -803 -219
rect -791 -219 -788 -201
rect -725 -206 -722 -191
rect -728 -211 -722 -206
rect -798 -222 -788 -219
<< m123contact >>
rect -790 303 -785 308
rect -623 303 -618 308
rect -516 291 -511 296
rect -403 291 -398 296
rect -203 291 -198 296
rect -97 291 -92 296
rect -801 275 -796 280
rect -788 279 -783 284
rect -766 276 -761 281
rect -742 272 -737 277
rect -671 272 -666 277
rect -659 272 -654 277
rect -647 276 -642 281
rect -625 279 -620 284
rect -612 275 -607 280
rect -814 248 -809 253
rect -763 255 -758 260
rect -650 255 -645 260
rect -787 241 -782 246
rect -775 234 -770 239
rect -564 260 -559 265
rect -552 260 -547 265
rect -540 264 -535 269
rect -518 267 -513 272
rect -505 263 -500 268
rect -414 263 -409 268
rect -401 267 -396 272
rect -379 264 -374 269
rect -599 248 -594 253
rect -638 234 -633 239
rect -543 243 -538 248
rect -367 260 -362 265
rect -355 260 -350 265
rect -251 260 -246 265
rect -239 260 -234 265
rect -227 264 -222 269
rect -205 267 -200 272
rect -192 263 -187 268
rect -145 260 -140 265
rect -133 260 -128 265
rect -121 264 -116 269
rect -99 267 -94 272
rect -86 263 -81 268
rect -492 236 -487 241
rect -531 222 -526 227
rect -427 236 -422 241
rect -376 243 -371 248
rect -230 243 -225 248
rect -388 222 -383 227
rect -124 243 -119 248
rect -179 236 -174 241
rect -218 222 -213 227
rect -73 236 -68 241
rect -112 222 -107 227
rect -778 208 -773 213
rect -705 208 -700 213
rect -640 202 -635 207
rect -720 193 -715 198
rect -648 193 -643 198
rect -788 185 -783 190
rect -759 158 -754 163
rect -750 185 -745 190
rect -678 185 -673 190
rect -713 158 -708 163
rect -687 158 -682 163
rect -750 122 -745 127
rect -678 122 -673 127
rect -781 92 -776 97
rect -698 92 -693 97
rect -802 40 -797 45
rect -779 39 -774 44
rect -758 39 -753 44
rect -749 39 -744 44
rect -737 39 -732 44
rect -728 39 -723 44
rect -716 39 -711 44
rect -707 39 -702 44
rect -695 39 -690 44
rect -869 -50 -864 -45
rect -652 113 -646 118
rect -2 218 3 223
rect -601 196 -596 201
rect -528 196 -523 201
rect -417 196 -412 201
rect -344 196 -339 201
rect -235 196 -230 201
rect -162 196 -157 201
rect -463 190 -458 195
rect -279 190 -274 195
rect -97 190 -92 195
rect -543 181 -538 186
rect -471 181 -466 186
rect -582 146 -577 151
rect -573 173 -568 178
rect -501 173 -496 178
rect -536 146 -531 151
rect -510 146 -505 151
rect -573 110 -568 115
rect -501 110 -496 115
rect -678 77 -673 82
rect -653 77 -648 82
rect -625 77 -620 82
rect -475 101 -469 106
rect -359 181 -354 186
rect -287 181 -282 186
rect -398 146 -393 151
rect -389 173 -384 178
rect -317 173 -312 178
rect -352 146 -347 151
rect -326 146 -321 151
rect -389 110 -384 115
rect -317 110 -312 115
rect -501 65 -496 70
rect -476 65 -471 70
rect -448 65 -443 70
rect -291 101 -285 106
rect -177 181 -172 186
rect -105 181 -100 186
rect -216 146 -211 151
rect -207 173 -202 178
rect -170 146 -165 151
rect -144 146 -139 151
rect -207 110 -202 115
rect -135 110 -130 115
rect -317 65 -312 70
rect -292 65 -287 70
rect -264 65 -259 70
rect -50 187 -45 192
rect -26 191 -21 196
rect -4 194 1 199
rect 9 190 14 195
rect -29 170 -24 175
rect 22 163 27 168
rect -5 156 0 161
rect -17 149 -12 154
rect -12 140 -7 145
rect -60 109 -55 114
rect -36 113 -31 118
rect -14 116 -9 121
rect -1 112 4 117
rect -109 101 -103 106
rect -39 92 -34 97
rect -54 73 -49 78
rect 12 85 17 90
rect -15 78 -10 83
rect -27 71 -22 76
rect -135 65 -130 70
rect -110 65 -105 70
rect -82 65 -77 70
rect -26 62 -21 67
rect -573 56 -568 61
rect -389 56 -384 61
rect -207 56 -202 61
rect -674 45 -669 50
rect -476 40 -471 45
rect -497 35 -492 40
rect -476 26 -471 31
rect -498 15 -493 20
rect -368 39 -363 44
rect -325 40 -320 45
rect -292 40 -287 45
rect -332 31 -327 36
rect -313 33 -308 38
rect -292 26 -287 31
rect -314 15 -309 20
rect -425 3 -420 8
rect -413 3 -408 8
rect -404 3 -399 8
rect -392 3 -387 8
rect -383 3 -378 8
rect -371 3 -366 8
rect -647 -5 -642 0
rect -635 -5 -630 0
rect -626 -5 -621 0
rect -614 -5 -609 0
rect -605 -5 -600 0
rect -593 -5 -588 0
rect -584 -5 -579 0
rect -562 -5 -557 0
rect -477 -3 -472 2
rect -655 -14 -650 -9
rect -705 -41 -700 -36
rect -684 -41 -679 -36
rect -668 -41 -663 -36
rect -846 -50 -841 -45
rect -828 -50 -823 -45
rect -816 -50 -811 -45
rect -807 -50 -802 -45
rect -795 -50 -790 -45
rect -786 -50 -781 -45
rect -774 -50 -769 -45
rect -765 -50 -760 -45
rect -721 -48 -716 -43
rect -853 -68 -848 -63
rect -748 -58 -743 -53
rect -749 -76 -744 -71
rect -667 -73 -662 -68
rect -508 -10 -503 -5
rect -448 -10 -443 -5
rect -547 -48 -542 -43
rect -575 -54 -570 -49
rect -575 -63 -570 -58
rect -783 -105 -778 -100
rect -644 -116 -639 -111
rect -632 -116 -627 -111
rect -623 -116 -618 -111
rect -611 -116 -606 -111
rect -602 -116 -597 -111
rect -590 -116 -585 -111
rect -469 -45 -464 -40
rect -437 -46 -432 -41
rect -508 -55 -503 -50
rect -488 -78 -483 -73
rect -424 -76 -419 -71
rect -559 -91 -554 -86
rect -547 -91 -542 -86
rect -538 -91 -533 -86
rect -526 -91 -521 -86
rect -517 -91 -512 -86
rect -505 -91 -500 -86
rect -439 -91 -434 -86
rect -293 6 -288 11
rect -110 44 -105 49
rect -131 35 -126 40
rect -213 26 -208 31
rect -110 26 -105 31
rect -241 21 -236 26
rect -132 15 -127 20
rect -332 -2 -327 3
rect -214 1 -209 6
rect -342 -11 -337 -6
rect -325 -11 -320 -6
rect -374 -36 -369 -31
rect -352 -43 -347 -38
rect -111 -3 -106 2
rect -178 -8 -173 -3
rect -143 -8 -138 -3
rect -285 -45 -280 -40
rect -262 -46 -257 -41
rect -213 -46 -208 -41
rect -103 -45 -98 -40
rect -71 -46 -66 -41
rect -37 34 -32 39
rect -24 38 -19 43
rect -2 35 3 40
rect 22 31 27 36
rect -50 7 -45 12
rect 1 14 6 19
rect -23 0 -18 5
rect -11 -7 -6 -2
rect 1 -25 6 -20
rect -325 -51 -320 -46
rect -253 -53 -248 -48
rect -47 -56 -42 -51
rect -35 -56 -30 -51
rect -23 -52 -18 -47
rect -1 -49 4 -44
rect 12 -53 17 -48
rect -304 -78 -299 -73
rect -375 -88 -370 -83
rect -363 -88 -358 -83
rect -354 -88 -349 -83
rect -567 -105 -562 -100
rect -737 -127 -732 -122
rect -725 -127 -720 -122
rect -716 -127 -711 -122
rect -704 -127 -699 -122
rect -695 -127 -690 -122
rect -683 -127 -678 -122
rect -674 -127 -669 -122
rect -662 -127 -657 -122
rect -782 -146 -777 -141
rect -818 -153 -813 -148
rect -829 -181 -824 -176
rect -816 -177 -811 -172
rect -794 -180 -789 -175
rect -569 -128 -564 -123
rect -342 -88 -337 -83
rect -333 -88 -328 -83
rect -321 -88 -316 -83
rect -264 -102 -259 -97
rect -170 -62 -165 -57
rect -26 -73 -21 -68
rect -199 -78 -194 -73
rect -122 -78 -117 -73
rect 25 -80 30 -75
rect -14 -94 -9 -89
rect -210 -106 -205 -101
rect -197 -102 -192 -97
rect -175 -105 -170 -100
rect -163 -109 -158 -104
rect -151 -109 -146 -104
rect -508 -130 -503 -125
rect -468 -127 -463 -122
rect -456 -127 -451 -122
rect -447 -127 -442 -122
rect -435 -127 -430 -122
rect -426 -127 -421 -122
rect -414 -127 -409 -122
rect -405 -127 -400 -122
rect -393 -127 -388 -122
rect -223 -133 -218 -128
rect -172 -126 -167 -121
rect -184 -147 -179 -142
rect -14 -103 -9 -98
rect -26 -124 -21 -119
rect 25 -117 30 -112
rect -47 -141 -42 -136
rect -35 -141 -30 -136
rect -23 -145 -18 -140
rect -1 -148 4 -143
rect 12 -144 17 -139
rect -616 -167 -611 -162
rect -396 -176 -391 -171
rect 1 -172 6 -167
rect -782 -184 -777 -179
rect -770 -184 -765 -179
rect -842 -208 -837 -203
rect -607 -189 -602 -184
rect -791 -201 -786 -196
rect -803 -222 -798 -217
<< metal3 >>
rect -785 303 -784 307
rect -787 284 -784 303
rect -624 303 -623 307
rect -624 284 -621 303
rect -517 291 -516 295
rect -398 291 -397 295
rect -517 272 -514 291
rect -400 272 -397 291
rect -204 291 -203 295
rect -98 291 -97 295
rect -204 272 -201 291
rect -98 272 -95 291
rect -681 226 -595 230
rect -773 208 -705 213
rect -778 114 -773 208
rect -681 198 -676 226
rect -598 218 -595 226
rect -3 218 -2 222
rect -598 215 0 218
rect -598 214 -315 215
rect -715 194 -648 198
rect -652 193 -648 194
rect -596 196 -528 201
rect -652 118 -646 193
rect -778 111 -682 114
rect -698 97 -695 111
rect -685 92 -682 111
rect -601 92 -596 196
rect -504 186 -499 214
rect -412 196 -344 201
rect -538 182 -471 186
rect -475 181 -471 182
rect -475 106 -469 181
rect -417 92 -412 196
rect -320 186 -315 214
rect -230 196 -162 201
rect -354 182 -287 186
rect -291 181 -287 182
rect -291 106 -285 181
rect -235 92 -230 196
rect -138 186 -133 215
rect -3 199 0 215
rect -172 182 -105 186
rect -109 181 -105 182
rect -109 144 -103 181
rect -109 141 -12 144
rect -109 106 -103 141
rect -13 140 -12 141
rect -13 121 -10 140
rect -685 89 -230 92
rect -685 50 -682 89
rect -685 46 -674 50
rect -811 41 -802 44
rect -811 -6 -808 41
rect -693 5 -690 39
rect -601 40 -596 89
rect -417 52 -412 89
rect -417 49 -310 52
rect -601 36 -497 40
rect -836 -9 -808 -6
rect -705 2 -690 5
rect -836 -56 -833 -9
rect -705 -36 -702 2
rect -683 -45 -680 -41
rect -716 -48 -680 -45
rect -756 -56 -748 -53
rect -836 -59 -766 -56
rect -769 -99 -766 -59
rect -769 -102 -760 -99
rect -763 -119 -760 -102
rect -756 -112 -753 -56
rect -665 -54 -575 -51
rect -570 -54 -567 36
rect -363 40 -325 44
rect -363 39 -347 40
rect -313 38 -310 49
rect -235 40 -230 89
rect -61 74 -54 77
rect -61 40 -58 74
rect -21 62 -20 66
rect -23 43 -20 62
rect -235 36 -131 40
rect -235 26 -230 36
rect -126 36 -58 40
rect -236 21 -230 26
rect -508 -50 -505 -10
rect -665 -68 -662 -54
rect -736 -71 -667 -68
rect -736 -72 -733 -71
rect -744 -75 -733 -72
rect -496 -73 -493 15
rect -496 -77 -488 -73
rect -756 -115 -644 -112
rect -763 -122 -741 -119
rect -813 -153 -812 -149
rect -815 -172 -812 -153
rect -744 -152 -741 -122
rect -496 -125 -493 -77
rect -446 -83 -443 -10
rect -435 -11 -342 -8
rect -435 -41 -432 -11
rect -313 -31 -309 15
rect -173 -7 -143 -3
rect -369 -34 -309 -31
rect -437 -58 -434 -46
rect -313 -73 -309 -34
rect -131 -12 -127 15
rect 55 9 60 14
rect -11 -11 -8 -7
rect 55 -11 58 9
rect -11 -12 58 -11
rect -131 -14 58 -12
rect -131 -15 -8 -14
rect -131 -73 -127 -15
rect 0 -25 1 -21
rect 0 -44 3 -25
rect -313 -77 -304 -73
rect -194 -78 -193 -74
rect -131 -77 -122 -73
rect -446 -86 -434 -83
rect -196 -97 -193 -78
rect -503 -128 -493 -125
rect -497 -132 -493 -128
rect -497 -135 -393 -132
rect -744 -155 -611 -152
rect -614 -162 -611 -155
rect -396 -171 -393 -135
rect 0 -167 3 -148
rect 0 -171 1 -167
rect -815 -193 -812 -177
rect -823 -196 -812 -193
rect -823 -226 -820 -196
rect -774 -226 -769 -225
rect -823 -229 -769 -226
rect -774 -230 -769 -229
<< m234contact >>
rect -806 63 -801 68
rect -653 63 -648 68
rect -660 -25 -655 -20
rect -659 -41 -654 -36
rect -524 -41 -519 -36
rect -486 -3 -481 2
rect -721 -81 -716 -76
rect -438 -63 -433 -58
rect -409 -60 -404 -55
rect -579 -137 -574 -132
rect -540 -152 -535 -147
<< metal4 >>
rect -801 64 -653 67
rect -667 12 -502 15
rect -667 -29 -664 12
rect -505 2 -502 12
rect -505 -1 -486 2
rect -655 -23 -531 -20
rect -667 -32 -656 -29
rect -659 -36 -656 -32
rect -650 -77 -647 -23
rect -534 -26 -531 -23
rect -534 -29 -521 -26
rect -524 -36 -521 -29
rect -408 -55 -405 -51
rect -437 -67 -434 -63
rect -716 -80 -647 -77
rect -578 -70 -434 -67
rect -578 -132 -575 -70
rect -408 -96 -405 -60
rect -539 -99 -405 -96
rect -539 -147 -536 -99
<< metal5 >>
rect -824 281 -95 284
rect -824 227 -821 281
rect -752 277 -749 281
rect -753 272 -748 277
rect -692 267 -687 272
rect -690 256 -687 267
rect -690 253 -674 256
rect -824 224 -802 227
rect -805 -112 -802 224
rect -677 150 -674 253
rect -624 246 -621 281
rect -583 251 -578 256
rect -625 241 -620 246
rect -581 222 -578 251
rect -517 234 -514 281
rect -478 266 -438 269
rect -518 229 -513 234
rect -616 219 -578 222
rect -678 145 -673 150
rect -625 149 -620 150
rect -616 149 -613 219
rect -609 177 -604 178
rect -478 177 -475 266
rect -443 264 -438 266
rect -272 259 -267 264
rect -165 259 -160 264
rect -272 258 -268 259
rect -609 174 -475 177
rect -463 255 -268 258
rect -609 173 -604 174
rect -625 146 -613 149
rect -625 145 -620 146
rect -501 135 -496 136
rect -463 135 -460 255
rect -163 247 -160 259
rect -447 244 -160 247
rect -447 148 -444 244
rect -98 234 -95 281
rect -401 233 -396 234
rect -205 233 -200 234
rect -99 233 -94 234
rect -401 230 -35 233
rect -401 229 -396 230
rect -205 229 -200 230
rect -99 229 -94 230
rect -38 192 -35 230
rect -75 186 -66 191
rect -39 190 -34 192
rect -43 187 -34 190
rect -427 173 -422 178
rect -245 173 -240 178
rect -135 176 -130 178
rect -75 176 -72 186
rect -135 173 -72 176
rect -43 174 -40 187
rect -448 143 -443 148
rect -426 142 -423 173
rect -264 147 -259 149
rect -264 144 -249 147
rect -426 139 -342 142
rect -501 132 -460 135
rect -501 131 -496 132
rect -345 -18 -342 139
rect -277 140 -272 141
rect -277 137 -256 140
rect -277 136 -272 137
rect -259 29 -256 137
rect -252 41 -249 144
rect -245 51 -242 173
rect -49 171 -40 174
rect -49 114 -46 171
rect -49 112 -44 114
rect 12 112 15 113
rect -49 109 15 112
rect -245 48 -68 51
rect -252 38 -84 41
rect -259 26 -97 29
rect -345 -21 -241 -18
rect -244 -100 -241 -21
rect -100 -80 -97 26
rect -87 18 -84 38
rect -71 31 -68 48
rect 12 44 15 109
rect 0 41 15 44
rect -59 31 -54 32
rect -71 28 -53 31
rect -59 27 -54 28
rect -87 15 -75 18
rect -78 -71 -75 15
rect -67 -65 -62 -60
rect -66 -71 -63 -65
rect -78 -74 -63 -71
rect -100 -83 -62 -80
rect 0 -82 3 41
rect 12 36 15 41
rect 11 31 16 36
rect 12 -25 17 -20
rect -237 -100 -232 -99
rect -244 -103 -232 -100
rect -237 -104 -232 -103
rect -844 -115 -802 -112
rect -844 -132 -841 -115
rect -783 -122 -778 -121
rect -829 -125 -778 -122
rect -829 -127 -824 -125
rect -783 -126 -778 -125
rect -65 -126 -62 -83
rect -1 -87 4 -82
rect 0 -95 3 -87
rect -40 -98 3 -95
rect -66 -131 -61 -126
rect -844 -135 -812 -132
rect -815 -210 -812 -135
rect -197 -136 -192 -135
rect -40 -136 -37 -98
rect 0 -105 3 -98
rect -1 -110 4 -105
rect -197 -139 -37 -136
rect -197 -140 -192 -139
rect 13 -168 16 -25
rect 12 -173 17 -168
rect -816 -215 -811 -210
<< pad >>
rect -753 272 -748 277
rect -692 267 -687 272
rect -443 264 -438 269
rect -272 259 -267 264
rect -165 259 -160 264
rect -583 251 -578 256
rect -625 241 -620 246
rect -518 229 -513 234
rect -401 229 -396 234
rect -205 229 -200 234
rect -99 229 -94 234
rect -71 186 -66 191
rect -39 187 -34 192
rect -609 173 -604 178
rect -427 173 -422 178
rect -245 173 -240 178
rect -135 173 -130 178
rect -678 145 -673 150
rect -625 145 -620 150
rect -448 143 -443 148
rect -264 144 -259 149
rect -277 136 -272 141
rect -501 131 -496 136
rect -49 109 -44 114
rect -59 27 -54 32
rect 11 31 16 36
rect 38 30 43 35
rect 53 30 58 35
rect 55 9 60 14
rect 12 -25 17 -20
rect -67 -65 -62 -60
rect -1 -87 4 -82
rect -237 -104 -232 -99
rect -130 -110 -125 -105
rect -1 -110 4 -105
rect -829 -127 -824 -122
rect -783 -126 -778 -121
rect -66 -131 -61 -126
rect -197 -140 -192 -135
rect -135 -156 -130 -151
rect 12 -173 17 -168
rect -755 -185 -750 -180
rect -816 -215 -811 -210
rect -728 -211 -723 -206
rect -774 -230 -769 -225
<< labels >>
rlabel metal3 -138 214 -133 218 1 vdd
rlabel m123contact -170 146 -165 151 1 p_0
rlabel metal1 -110 1 -106 5 1 g_0
rlabel m123contact -135 110 -130 115 1 b_0
rlabel metal2 -82 143 -77 148 1 a_0
rlabel m123contact -207 110 -202 115 1 c0
rlabel metal3 -235 36 -230 40 1 gnd
rlabel m123contact -352 146 -347 151 1 p_1
rlabel m123contact -389 110 -384 115 1 c1
rlabel m123contact -317 110 -312 115 1 b_1
rlabel metal1 -102 -44 -97 -41 1 p0c0
rlabel m123contact -292 26 -287 31 1 gb_1
rlabel m123contact -110 26 -105 31 1 gb_0
rlabel metal1 -284 -44 -279 -41 1 p1g0
rlabel m123contact -375 -88 -370 -83 1 p1p0c0
rlabel m123contact -573 110 -568 115 1 c2
rlabel metal2 -448 143 -443 148 1 a_2
rlabel m123contact -501 110 -496 115 1 b_2
rlabel m123contact -536 146 -531 151 1 p_2
rlabel metal1 -476 1 -472 5 1 g_2
rlabel m123contact -476 26 -471 31 1 gb_2
rlabel metal1 -468 -44 -463 -41 1 p2g1
rlabel m123contact -559 -91 -554 -86 1 p2p1g0
rlabel metal3 -468 -127 -463 -122 1 p2p1p0c0
rlabel metal2 -625 145 -620 150 1 a_3
rlabel m123contact -678 122 -673 127 1 b_3
rlabel m123contact -788 185 -783 190 3 s3
rlabel m123contact -293 6 -288 11 1 g_1
rlabel m123contact -697 94 -695 95 1 gnd
rlabel metal1 -668 -72 -664 -70 8 gnd
rlabel m123contact -704 -40 -701 -37 1 p_3
rlabel metal1 -688 -40 -684 -38 1 p3g2
rlabel metal1 -555 -53 -552 -52 1 vdd
rlabel metal1 -686 -5 -686 -5 1 vdd
rlabel metal1 -590 -157 -586 -156 8 gnd
rlabel m123contact -567 -105 -562 -100 1 p_2
rlabel metal1 -620 -79 -619 -78 1 vdd
rlabel polycontact -594 -115 -590 -111 1 p_3
rlabel m123contact -644 -116 -639 -111 1 p3p2g1
rlabel metal1 -689 -89 -685 -88 5 vdd
rlabel polycontact -687 -126 -683 -122 1 p_2
rlabel polycontact -708 -126 -704 -122 1 p_1
rlabel polycontact -530 -90 -526 -86 1 g_0
rlabel m123contact -737 -127 -732 -122 1 p3p2p1g0
rlabel metal1 -783 6 -783 6 1 vdd
rlabel metal1 -787 -12 -787 -12 1 vdd
rlabel metal1 -753 -96 -753 -96 1 gnd
rlabel metal1 -796 41 -796 41 1 p
rlabel metal1 -638 -171 -636 -167 4 gnd
rlabel metal1 -606 -191 -604 -187 3 out
rlabel metal1 -570 -180 -570 -180 1 vdd
rlabel metal1 -607 -170 -603 -165 1 p
rlabel metal1 -749 -107 -747 -103 6 gnd
rlabel metal1 -815 -131 -813 -118 3 vdd
rlabel metal1 -606 -210 -603 -204 1 c0
rlabel metal1 -781 -129 -779 -127 1 c4
rlabel m123contact -647 -5 -642 0 1 c3
rlabel m123contact -562 -5 -557 0 1 gb_2
rlabel m123contact -713 158 -708 163 1 p_3
rlabel m123contact -652 79 -652 79 1 gb_3
rlabel metal1 -866 -10 -866 -10 4 vdd
rlabel m123contact -781 -103 -781 -103 1 gb
rlabel m123contact -828 -50 -823 -45 1 g
rlabel metal1 1 138 4 141 5 vdd
rlabel metal2 14 72 17 74 1 gnd
rlabel metal1 -63 134 -60 137 5 vdd
rlabel metal1 -62 97 -59 99 1 gnd
rlabel m123contact -12 140 -7 145 5 vdd
rlabel metal1 -76 109 -73 113 1 a_0
rlabel metal1 20 113 23 116 1 a0_in
rlabel metal1 11 216 14 219 5 vdd
rlabel metal2 24 150 27 152 1 gnd
rlabel metal1 -53 212 -50 215 5 vdd
rlabel metal1 -52 175 -49 177 1 gnd
rlabel m123contact -17 149 -12 154 1 gnd
rlabel m123contact -2 218 3 223 5 vdd
rlabel metal1 -66 187 -63 191 1 b_0
rlabel metal1 30 191 33 194 1 b0_in
rlabel m123contact -27 71 -22 76 1 gnd
rlabel m123contact -26 62 -21 67 5 vdd
rlabel m123contact -11 -7 -6 -2 1 gnd
rlabel metal1 26 19 29 21 1 gnd
rlabel metal1 27 56 30 59 5 vdd
rlabel metal2 -50 -6 -47 -4 1 gnd
rlabel metal1 -37 60 -34 63 5 vdd
rlabel pad -245 173 -240 178 1 s0
rlabel pad -57 29 -55 30 1 s0
rlabel metal1 40 31 43 35 1 s0_out
rlabel polycontact 20 -141 24 -137 5 clk
rlabel metal1 14 -168 17 -165 1 vdd
rlabel metal2 27 -101 30 -99 5 gnd
rlabel polycontact -6 -165 -2 -161 1 clk
rlabel polycontact -6 -110 -2 -106 5 clk
rlabel polycontact -30 -140 -26 -136 5 clk
rlabel metal1 -50 -164 -47 -161 1 vdd
rlabel metal1 -49 -126 -46 -124 5 gnd
rlabel m123contact -14 -103 -9 -98 5 gnd
rlabel m123contact 1 -172 6 -167 1 vdd
rlabel polycontact 20 -55 24 -51 1 clk
rlabel metal1 14 -27 17 -24 5 vdd
rlabel metal2 27 -93 30 -91 1 gnd
rlabel polycontact -6 -31 -2 -27 5 clk
rlabel polycontact -6 -86 -2 -82 1 clk
rlabel polycontact -30 -56 -26 -52 1 clk
rlabel metal1 -50 -31 -47 -28 5 vdd
rlabel metal1 -49 -68 -46 -66 1 gnd
rlabel m123contact -14 -94 -9 -89 1 gnd
rlabel m123contact 1 -25 6 -20 5 vdd
rlabel metal1 33 -52 36 -49 1 a1_in
rlabel metal1 -63 -56 -60 -52 1 a_1
rlabel metal1 33 -143 36 -140 1 b1_in
rlabel polycontact -217 -108 -213 -104 1 clk
rlabel metal1 -210 -80 -207 -77 5 vdd
rlabel metal2 -223 -146 -220 -144 1 gnd
rlabel polycontact -191 -84 -187 -80 5 clk
rlabel polycontact -191 -139 -187 -135 1 clk
rlabel polycontact -167 -109 -163 -105 1 clk
rlabel metal1 -146 -84 -143 -81 5 vdd
rlabel metal1 -147 -121 -144 -119 1 gnd
rlabel m123contact -184 -147 -179 -142 1 gnd
rlabel m123contact -199 -78 -194 -73 5 vdd
rlabel metal1 -63 -140 -60 -136 1 b_1
rlabel pad -427 173 -422 178 1 s1
rlabel metal1 -229 -105 -226 -102 1 s1
rlabel metal1 -135 -109 -130 -105 1 s1_out
rlabel polycontact 6 31 10 35 1 clk
rlabel polycontact -18 56 -14 60 5 clk
rlabel polycontact -44 32 -40 36 1 clk
rlabel polycontact -18 1 -14 5 1 clk
rlabel polycontact -43 109 -39 113 1 clk
rlabel polycontact -19 134 -15 138 5 clk
rlabel polycontact 7 110 11 114 1 clk
rlabel polycontact -19 79 -15 83 1 clk
rlabel polycontact -33 187 -29 191 1 clk
rlabel polycontact -9 212 -5 216 5 clk
rlabel polycontact 17 188 21 192 1 clk
rlabel polycontact -9 157 -5 161 1 clk
rlabel metal2 -264 144 -259 149 1 a_1
rlabel polycontact -78 261 -74 265 1 clk
rlabel metal1 -84 289 -81 292 5 vdd
rlabel metal2 -71 223 -68 225 1 gnd
rlabel polycontact -104 285 -100 289 5 clk
rlabel polycontact -104 230 -100 234 1 clk
rlabel polycontact -128 260 -124 264 1 clk
rlabel metal1 -148 285 -145 288 5 vdd
rlabel metal1 -147 248 -144 250 1 gnd
rlabel m123contact -112 222 -107 227 1 gnd
rlabel m123contact -97 291 -92 296 5 vdd
rlabel polycontact -184 261 -180 265 1 clk
rlabel metal1 -190 289 -187 292 5 vdd
rlabel metal2 -177 223 -174 225 1 gnd
rlabel polycontact -210 285 -206 289 5 clk
rlabel polycontact -210 230 -206 234 1 clk
rlabel polycontact -234 260 -230 264 1 clk
rlabel metal1 -254 285 -251 288 5 vdd
rlabel metal1 -253 248 -250 250 1 gnd
rlabel m123contact -218 222 -213 227 1 gnd
rlabel m123contact -203 291 -198 296 5 vdd
rlabel metal1 -157 262 -157 262 1 a_2
rlabel metal1 -65 264 -62 267 1 a2_in
rlabel metal1 -267 260 -264 264 1 b_2
rlabel metal1 -171 264 -168 267 1 b2_in
rlabel polycontact -421 261 -417 265 1 clk
rlabel metal1 -414 289 -411 292 5 vdd
rlabel metal2 -427 223 -424 225 1 gnd
rlabel polycontact -395 285 -391 289 5 clk
rlabel polycontact -395 230 -391 234 1 clk
rlabel polycontact -371 260 -367 264 1 clk
rlabel metal1 -350 285 -347 288 5 vdd
rlabel metal1 -351 248 -348 250 1 gnd
rlabel m123contact -388 222 -383 227 1 gnd
rlabel m123contact -403 291 -398 296 5 vdd
rlabel pad -441 266 -441 266 1 s2
rlabel metal1 -337 260 -334 264 1 s2_out
rlabel polycontact -497 261 -493 265 1 clk
rlabel metal1 -503 289 -500 292 5 vdd
rlabel metal2 -490 223 -487 225 1 gnd
rlabel polycontact -523 285 -519 289 5 clk
rlabel polycontact -523 230 -519 234 1 clk
rlabel polycontact -547 260 -543 264 1 clk
rlabel metal1 -567 285 -564 288 5 vdd
rlabel metal1 -566 248 -563 250 1 gnd
rlabel m123contact -531 222 -526 227 1 gnd
rlabel m123contact -516 291 -511 296 5 vdd
rlabel polycontact -604 273 -600 277 1 clk
rlabel metal1 -610 301 -607 304 5 vdd
rlabel metal2 -597 235 -594 237 1 gnd
rlabel polycontact -630 297 -626 301 5 clk
rlabel polycontact -630 242 -626 246 1 clk
rlabel polycontact -654 272 -650 276 1 clk
rlabel metal1 -674 297 -671 300 5 vdd
rlabel metal1 -673 260 -670 262 1 gnd
rlabel m123contact -638 234 -633 239 1 gnd
rlabel m123contact -623 303 -618 308 5 vdd
rlabel pad -609 173 -604 178 1 s2
rlabel metal1 -580 260 -577 264 1 a_3
rlabel metal1 -484 264 -481 267 1 a3_in
rlabel metal1 -591 276 -588 279 1 b3_in
rlabel m123contact -818 -153 -813 -148 5 vdd
rlabel m123contact -803 -222 -798 -217 1 gnd
rlabel metal1 -766 -196 -763 -194 1 gnd
rlabel metal1 -765 -159 -762 -156 5 vdd
rlabel polycontact -786 -184 -782 -180 1 clk
rlabel polycontact -810 -214 -806 -210 1 clk
rlabel polycontact -810 -159 -806 -155 5 clk
rlabel metal2 -842 -221 -839 -219 1 gnd
rlabel metal1 -829 -155 -826 -152 5 vdd
rlabel polycontact -836 -183 -832 -179 1 clk
rlabel metal1 -848 -180 -845 -177 1 c4
rlabel metal1 -687 272 -684 276 1 b_3
rlabel metal1 -707 -231 -707 -231 8 gnd
rlabel metal1 -765 -231 -765 -231 2 vdd
rlabel metal1 -753 -184 -750 -180 1 c4_out
rlabel metal1 -730 -232 -726 -228 1 load1
rlabel metal1 -95 -177 -95 -177 8 vdd
rlabel metal1 -153 -177 -153 -177 2 gnd
rlabel metal1 -134 -178 -130 -175 1 load2
rlabel metal1 78 70 78 70 6 vdd
rlabel metal1 78 12 78 12 8 gnd
rlabel metal1 75 31 79 35 7 load3
rlabel metal1 -299 288 -299 288 6 vdd
rlabel metal1 -299 230 -299 230 8 gnd
rlabel metal1 -303 249 -298 253 1 load4
rlabel metal1 -724 272 -721 276 1 s3_out
rlabel metal1 -820 276 -817 279 1 s3
rlabel m123contact -790 303 -785 308 5 vdd
rlabel m123contact -775 234 -770 239 1 gnd
rlabel metal1 -738 260 -735 262 1 gnd
rlabel metal1 -737 297 -734 300 5 vdd
rlabel polycontact -758 272 -754 276 1 clk
rlabel polycontact -782 242 -778 246 1 clk
rlabel polycontact -782 297 -778 301 5 clk
rlabel metal2 -814 235 -811 237 1 gnd
rlabel metal1 -801 301 -798 304 5 vdd
rlabel polycontact -808 273 -804 277 1 clk
rlabel metal1 -696 299 -696 299 6 vdd
rlabel metal1 -696 241 -696 241 8 gnd
rlabel metal1 -701 260 -695 264 1 load5
<< end >>
