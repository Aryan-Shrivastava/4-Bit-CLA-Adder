.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'

va a gnd pulse 0 1.8 0ns 1ns 1ns 10ns 20ns
vb b gnd pulse 0 1.8 0ns 1ns 1ns 5ns 10ns
vc c gnd pulse 0 1.8 0ns 1ns 1ns 15ns 30ns

*******************************************************************************************************************************************************
* Nand Gate 3 input
.subckt nand_3_in y a b c vdd gnd 
    .param n={3}
    M1 y a vdd vdd CMOSP W={width_P} L={2*LAMBDA} AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
    M2 y b vdd vdd CMOSP W={width_P} L={2*LAMBDA} AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
    M3 y c vdd vdd CMOSP W={width_P} L={2*LAMBDA} AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}

    M4 y a t1 t1 CMOSN W={n*width_N} L={2*LAMBDA} AS={5*n*width_N*LAMBDA} PS={10*LAMBDA+2*n*width_N} AD={5*n*width_N*LAMBDA} PD={10*LAMBDA+2*n*width_N}
    M5 t1 b t2 t2 CMOSN W={n*width_N} L={2*LAMBDA} AS={5*n*width_N*LAMBDA} PS={10*LAMBDA+2*n*width_N} AD={5*n*width_N*LAMBDA} PD={10*LAMBDA+2*n*width_N}
    M6 t2 c gnd gnd CMOSN W={n*width_N} L={2*LAMBDA} AS={5*n*width_N*LAMBDA} PS={10*LAMBDA+2*n*width_N} AD={5*n*width_N*LAMBDA} PD={10*LAMBDA+2*n*width_N}
.ends nand_3_in

x_nand_3_in y a b c vdd gnd nand_3_in

.tran 0.1n 100n
.control
    run
    set curplottitle="2023102025- Aryan Shrivastava"
    set color0=white
    set color1=black
    plot v(a) v(b)+2 v(c)+4 v(y)+6
.endc