.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'

va a gnd pulse 0 1.8 0ns 1ns 1ns 10ns 20ns
vb b gnd pulse 0 1.8 0ns 1ns 1ns 5ns 10ns

.option scale=0.09u



* SPICE3 file created from xor.ext - technology: scmos

.option scale=0.09u

M1000 a_bar a vdd w_n30_42# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 out b a_bar Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=100 ps=60
M1002 out a_bar b Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1003 a_bar a gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=50 ps=30
M1004 b a out w_30_50# CMOSP w=20 l=2
+  ad=100 pd=50 as=200 ps=100
M1005 out b a w_0_49# CMOSP w=20 l=2
+  ad=0 pd=0 as=100 ps=50
C0 a vdd 0.38fF
C1 b w_0_49# 0.07fF
C2 a_bar out 0.20fF
C3 a w_0_49# 0.09fF
C4 w_30_50# b 0.09fF
C5 w_30_50# a 0.07fF
C6 a_bar vdd 0.25fF
C7 a w_n30_42# 0.07fF
C8 a_bar w_n30_42# 0.05fF
C9 out w_0_49# 0.05fF
C10 a_bar b 0.11fF
C11 a a_bar 0.05fF
C12 a gnd 0.05fF
C13 w_30_50# out 0.05fF
C14 b out 0.63fF
C15 a out 0.38fF
C16 a_bar gnd 0.10fF
C17 vdd w_n30_42# 0.09fF
C18 gnd Gnd 0.03fF
C19 out Gnd 0.20fF
C20 a_bar Gnd 0.41fF
C21 vdd Gnd 0.03fF
C22 a Gnd 0.28fF
C23 b Gnd 0.84fF
C24 w_30_50# Gnd 0.80fF
C25 w_0_49# Gnd 0.67fF
C26 w_n30_42# Gnd 0.84fF

.tran 0.1n 50ns

.control
run
set color0=white
set color1=black
set curplottitle="2023102025- Aryan Shrivastava"
plot v(a) v(b)+2 v(out)+4
.endc
