magic
tech scmos
timestamp 1731414890
<< nwell >>
rect -44 29 0 63
<< ntransistor >>
rect -33 1 -31 21
rect -13 1 -11 21
<< ptransistor >>
rect -33 35 -31 55
rect -13 35 -11 55
<< ndiffusion >>
rect -34 1 -33 21
rect -31 1 -30 21
rect -14 1 -13 21
rect -11 1 -10 21
<< pdiffusion >>
rect -34 35 -33 55
rect -31 35 -30 55
rect -14 35 -13 55
rect -11 35 -10 55
<< ndcontact >>
rect -38 1 -34 21
rect -30 1 -26 21
rect -18 1 -14 21
rect -10 1 -6 21
<< pdcontact >>
rect -38 35 -34 55
rect -30 35 -26 55
rect -18 35 -14 55
rect -10 35 -6 55
<< polysilicon >>
rect -33 55 -31 58
rect -13 55 -11 58
rect -33 21 -31 35
rect -13 21 -11 35
rect -33 -3 -31 1
rect -13 -3 -11 1
<< polycontact >>
rect -37 24 -33 28
rect -11 24 -7 28
<< metal1 >>
rect -44 59 0 63
rect -38 55 -34 59
rect -10 55 -6 59
rect -30 28 -26 35
rect -18 28 -14 35
rect -44 24 -37 28
rect -30 25 -14 28
rect -18 21 -14 25
rect -7 24 0 28
rect -38 -4 -34 1
rect -30 -4 -26 1
rect -10 -4 -6 1
rect -42 -8 -33 -4
rect -30 -8 -6 -4
<< labels >>
rlabel metal1 -26 59 -13 61 5 vdd
rlabel metal1 -43 25 -39 27 3 a
rlabel metal1 -21 25 -17 27 1 out
rlabel metal1 -41 -7 -37 -5 2 gnd
rlabel metal1 -5 25 -1 27 7 b
<< end >>
