.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
va in gnd pulse (0 1.8 0 0.1n 0.1n 1n 2n)
* SPICE3 file created from inverter.ext - technology: scmos

.option scale=0.09u

M1000 out in vdd w_39_19# CMOSP w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 out in gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=50 ps=30
C0 w_39_19# vdd 0.09fF
C1 in gnd 0.05fF
C2 in out 0.05fF
C3 out w_39_19# 0.05fF
C4 in w_39_19# 0.07fF
C5 out vdd 0.25fF
C6 out gnd 0.14fF
C7 gnd Gnd 0.08fF
C8 out Gnd 0.06fF
C9 vdd Gnd 0.03fF
C10 in Gnd 0.13fF
C11 w_39_19# Gnd 0.84fF
.tran 0.1n 20n

.control
set color0=white
run 
plot v(in) v(out)+2
.endc