magic
tech scmos
timestamp 1732080899
<< nwell >>
rect -14 -11 85 12
rect -14 -34 10 -11
<< ntransistor >>
rect 23 -24 25 -19
rect 47 -24 49 -19
rect 71 -24 73 -19
rect 23 -39 25 -34
rect 47 -38 49 -33
rect -3 -45 -1 -40
<< ptransistor >>
rect -3 -4 -1 6
rect 23 -4 25 6
rect 47 -4 49 6
rect 71 -5 73 5
rect -3 -28 -1 -18
<< ndiffusion >>
rect 22 -24 23 -19
rect 25 -24 26 -19
rect 46 -24 47 -19
rect 49 -24 50 -19
rect 70 -24 71 -19
rect 73 -24 74 -19
rect 22 -39 23 -34
rect 25 -39 26 -34
rect 46 -38 47 -33
rect 49 -38 50 -33
rect -4 -45 -3 -40
rect -1 -45 0 -40
<< pdiffusion >>
rect -4 -4 -3 6
rect -1 -4 0 6
rect 22 -4 23 6
rect 25 -4 26 6
rect 46 -4 47 6
rect 49 -4 50 6
rect 70 -5 71 5
rect 73 -5 74 5
rect -4 -28 -3 -18
rect -1 -28 0 -18
<< ndcontact >>
rect 18 -24 22 -19
rect 26 -24 30 -19
rect 42 -24 46 -19
rect 50 -24 54 -19
rect 66 -24 70 -19
rect 74 -24 78 -19
rect 18 -39 22 -34
rect 26 -39 30 -34
rect 42 -38 46 -33
rect 50 -38 54 -33
rect -8 -45 -4 -40
rect 0 -45 4 -40
<< pdcontact >>
rect -8 -4 -4 6
rect 0 -4 4 6
rect 18 -4 22 6
rect 26 -4 30 6
rect 42 -4 46 6
rect 50 -4 54 6
rect 66 -5 70 5
rect 74 -5 78 5
rect -8 -28 -4 -18
rect 0 -28 4 -18
<< polysilicon >>
rect -3 6 -1 9
rect 23 6 25 9
rect 47 6 49 9
rect 71 5 73 8
rect -3 -7 -1 -4
rect 23 -7 25 -4
rect 47 -7 49 -4
rect -3 -18 -1 -15
rect 23 -19 25 -16
rect 47 -19 49 -16
rect 71 -19 73 -5
rect 23 -27 25 -24
rect 47 -27 49 -24
rect 71 -27 73 -24
rect -3 -31 -1 -28
rect 23 -34 25 -31
rect 47 -33 49 -30
rect -3 -40 -1 -37
rect 23 -42 25 -39
rect 47 -41 49 -38
rect -3 -48 -1 -45
<< polycontact >>
rect -4 9 0 13
rect 22 9 26 13
rect 46 9 50 13
rect -4 -15 0 -11
rect 22 -16 26 -12
rect 46 -16 50 -12
rect 67 -16 71 -12
rect 22 -46 26 -42
rect 46 -45 50 -41
rect -4 -52 0 -48
<< metal1 >>
rect 3 16 14 19
rect -16 9 -4 12
rect -16 -48 -13 9
rect 3 6 6 16
rect 19 16 70 19
rect -10 -4 -8 -1
rect 4 3 6 6
rect 9 9 22 12
rect 33 9 46 12
rect -10 -18 -7 -4
rect 9 -7 12 9
rect 33 -1 36 9
rect 53 6 56 16
rect 30 -4 36 -1
rect 40 -4 42 -1
rect 54 3 56 6
rect 66 5 70 16
rect 6 -8 12 -7
rect -3 -11 3 -9
rect 0 -12 3 -11
rect 8 -10 12 -8
rect 8 -12 9 -10
rect 12 -16 22 -13
rect -10 -21 -8 -18
rect 12 -21 15 -16
rect 29 -19 32 -4
rect 40 -7 43 -4
rect 4 -24 15 -21
rect 30 -21 32 -19
rect 40 -19 43 -12
rect 74 -12 78 -5
rect 74 -16 83 -12
rect 74 -19 78 -16
rect 1 -40 4 -28
rect 18 -34 21 -24
rect 30 -25 33 -21
rect 40 -22 42 -19
rect 54 -24 55 -21
rect 30 -28 38 -25
rect 30 -39 32 -36
rect -16 -51 -4 -48
rect 29 -49 32 -39
rect 35 -41 38 -28
rect 52 -33 55 -24
rect 66 -25 70 -24
rect 54 -36 55 -33
rect 58 -28 70 -25
rect 35 -44 46 -41
rect 58 -51 61 -28
rect 34 -54 61 -51
<< metal2 >>
rect 40 -7 65 -4
rect 62 -11 65 -7
rect 5 -16 8 -13
rect 5 -19 55 -16
rect -10 -51 -7 -40
rect 5 -42 8 -19
rect 5 -45 17 -42
rect -10 -54 29 -51
rect 41 -51 44 -33
rect 34 -54 44 -51
<< m123contact >>
rect 14 15 19 20
rect 3 -13 8 -8
rect 16 -9 21 -4
rect 38 -12 43 -7
rect 50 -16 55 -11
rect 62 -16 67 -11
rect -10 -40 -5 -35
rect 41 -33 46 -28
rect 17 -47 22 -42
rect 29 -54 34 -49
<< metal3 >>
rect 19 15 20 19
rect 17 -4 20 15
<< labels >>
rlabel metal1 -16 -12 -13 -9 3 d
rlabel polycontact -4 -15 0 -11 1 clk
rlabel metal1 3 13 6 16 5 vdd
rlabel metal2 -10 -53 -7 -51 1 gnd
rlabel polycontact 22 9 26 13 5 clk
rlabel polycontact 22 -46 26 -42 1 clk
rlabel polycontact 46 -16 50 -12 1 clk
rlabel metal1 67 9 70 12 5 vdd
rlabel metal1 66 -28 69 -26 1 gnd
rlabel metal1 80 -16 83 -12 1 q
rlabel m123contact 29 -54 34 -49 1 gnd
rlabel m123contact 14 15 19 20 5 vdd
<< end >>
