.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.param wp={10*LAMBDA}
.param wn={5*LAMBDA}
.global gnd vdd
Vdd	vdd	gnd	'SUPPLY'
va a gnd pulse  0 1.8 0ns 0ns 0ns 8ns 16ns
vclk clk gnd pulse 0 1.8 0ns 0ns 0ns 5ns 10ns

*******************************************************************************************************************************************************
* Inverter Circuit
.subckt inv y x vdd gnd 
    M1 y x gnd gnd  CMOSN W={width_N} L={2*LAMBDA} AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    M2 y x vdd vdd  CMOSP W={width_P} L={2*LAMBDA} AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv


*************************************************************************************************************************************************
.subckt flop out in clk vdd gnd
    *First Stage
    Mp3 temp1 in vdd vdd CMOSP L={2*LAMBDA} W={wp} AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
    Mp2 out_int1 clk temp1 vdd CMOSP L={2*LAMBDA} W={wp} AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
    Mn1 out_int1 in gnd gnd CMOSN L={2*LAMBDA} W={wn} AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
    *Second Stage
    Mp6 out_int2 clk vdd vdd CMOSP L={2*LAMBDA} W={wp} AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
    Mn5 out_int2 out_int1 temp2 gnd CMOSN L={2*LAMBDA} W={wn} AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
    Mn4 temp2 clk gnd gnd CMOSN L={2*LAMBDA} W={wn} AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn} 
    *Third Stage
    Mp9 out_int3 out_int2 vdd vdd CMOSP L={2*LAMBDA} W={wp} AS={5*wp*LAMBDA} PS={10*LAMBDA+2*wp} AD={5*wp*LAMBDA} PD={10*LAMBDA+2*wp}
    Mn8 out_int3 clk temp3 gnd CMOSN L={2*LAMBDA} W={wn} AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
    Mn7 temp3 out_int2 gnd gnd CMOSN L={2*LAMBDA} W={wn} AS={5*wn*LAMBDA} PS={10*LAMBDA+2*wn} AD={5*wn*LAMBDA} PD={10*LAMBDA+2*wn}
    *Inverter
    xinv out out_int3 vdd gnd inv
.ends flop

x_ff out a clk vdd gnd flop

.ic v(out)=0
.tran 0.001n 30n
.measure tran TPCQ TRIG v(clk) VAL='SUPPLY/2' RISE=3 TARG v(out) VAL='SUPPLY/2' RISE=2
.control
    run
    set curplottitle="2023102025- Aryan Shrivastava"
    set color0=white
    set color1=black
    plot v(a)+2 v(out)+4 v(clk)
.endc