magic
tech scmos
timestamp 1731596994
<< nwell >>
rect -751 194 -716 218
rect -682 194 -644 218
rect -744 164 -708 188
rect -672 164 -636 188
rect -574 182 -539 206
rect -505 182 -467 206
rect -390 182 -355 206
rect -321 182 -283 206
rect -208 182 -173 206
rect -139 182 -101 206
rect -743 123 -719 158
rect -671 123 -647 158
rect -567 152 -531 176
rect -495 152 -459 176
rect -383 152 -347 176
rect -311 152 -275 176
rect -201 152 -165 176
rect -129 152 -93 176
rect -676 83 -652 117
rect -646 83 -622 117
rect -566 111 -542 146
rect -494 111 -470 146
rect -382 111 -358 146
rect -310 111 -286 146
rect -200 111 -176 146
rect -128 111 -104 146
rect -499 71 -475 105
rect -469 71 -445 105
rect -315 71 -291 105
rect -285 71 -261 105
rect -133 71 -109 105
rect -103 71 -79 105
rect -800 4 -688 38
rect -652 1 -565 35
rect -471 1 -436 25
rect -430 9 -364 43
rect -287 1 -252 25
rect -867 -44 -843 -9
rect -833 -44 -746 -10
rect -705 -36 -661 -2
rect -487 -40 -443 -6
rect -303 -40 -259 -6
rect -208 -13 -174 31
rect -105 1 -70 25
rect -121 -40 -77 -6
rect -817 -144 -783 -100
rect -742 -121 -655 -87
rect -649 -110 -583 -76
rect -564 -85 -498 -51
rect -380 -82 -314 -48
rect -473 -121 -386 -87
rect -602 -210 -568 -164
<< ntransistor >>
rect -769 205 -759 207
rect -700 205 -690 207
rect -592 193 -582 195
rect -523 193 -513 195
rect -408 193 -398 195
rect -339 193 -329 195
rect -226 193 -216 195
rect -157 193 -147 195
rect -762 175 -752 177
rect -693 175 -683 177
rect -585 163 -575 165
rect -516 163 -506 165
rect -401 163 -391 165
rect -332 163 -322 165
rect -219 163 -209 165
rect -150 163 -140 165
rect -758 131 -756 141
rect -689 131 -687 141
rect -581 119 -579 129
rect -512 119 -510 129
rect -397 119 -395 129
rect -328 119 -326 129
rect -215 119 -213 129
rect -146 119 -144 129
rect -789 46 -787 56
rect -764 47 -762 87
rect -743 47 -741 87
rect -722 47 -720 87
rect -701 47 -699 87
rect -665 55 -663 75
rect -635 55 -633 75
rect -488 43 -486 63
rect -458 43 -456 63
rect -304 43 -302 63
rect -274 43 -272 63
rect -122 43 -120 63
rect -92 43 -90 63
rect -489 12 -479 14
rect -236 18 -216 20
rect -305 12 -295 14
rect -123 12 -113 14
rect -856 -62 -854 -52
rect -822 -93 -820 -53
rect -801 -93 -799 -53
rect -780 -93 -778 -53
rect -759 -93 -757 -53
rect -694 -64 -692 -44
rect -674 -64 -672 -44
rect -641 -48 -639 -8
rect -620 -48 -618 -8
rect -599 -48 -597 -8
rect -578 -48 -576 -8
rect -419 -30 -417 0
rect -398 -30 -396 0
rect -377 -30 -375 0
rect -236 -2 -216 0
rect -476 -68 -474 -48
rect -456 -68 -454 -48
rect -292 -68 -290 -48
rect -272 -68 -270 -48
rect -110 -68 -108 -48
rect -90 -68 -88 -48
rect -775 -113 -755 -111
rect -775 -133 -755 -131
rect -731 -170 -729 -130
rect -710 -170 -708 -130
rect -689 -170 -687 -130
rect -668 -170 -666 -130
rect -638 -149 -636 -119
rect -617 -149 -615 -119
rect -596 -149 -594 -119
rect -553 -124 -551 -94
rect -532 -124 -530 -94
rect -511 -124 -509 -94
rect -369 -121 -367 -91
rect -348 -121 -346 -91
rect -327 -121 -325 -91
rect -462 -170 -460 -130
rect -441 -170 -439 -130
rect -420 -170 -418 -130
rect -399 -170 -397 -130
rect -630 -177 -610 -175
rect -630 -199 -610 -197
<< ptransistor >>
rect -744 205 -724 207
rect -672 205 -652 207
rect -567 193 -547 195
rect -495 193 -475 195
rect -383 193 -363 195
rect -311 193 -291 195
rect -201 193 -181 195
rect -129 193 -109 195
rect -737 175 -717 177
rect -665 175 -645 177
rect -560 163 -540 165
rect -488 163 -468 165
rect -376 163 -356 165
rect -304 163 -284 165
rect -194 163 -174 165
rect -122 163 -102 165
rect -732 131 -730 151
rect -660 131 -658 151
rect -555 119 -553 139
rect -483 119 -481 139
rect -371 119 -369 139
rect -299 119 -297 139
rect -189 119 -187 139
rect -117 119 -115 139
rect -665 89 -663 109
rect -635 89 -633 109
rect -488 77 -486 97
rect -458 77 -456 97
rect -304 77 -302 97
rect -274 77 -272 97
rect -122 77 -120 97
rect -92 77 -90 97
rect -789 12 -787 32
rect -764 12 -762 32
rect -743 12 -741 32
rect -722 12 -720 32
rect -701 12 -699 32
rect -641 7 -639 27
rect -620 7 -618 27
rect -599 7 -597 27
rect -578 7 -576 27
rect -419 15 -417 35
rect -398 15 -396 35
rect -377 15 -375 35
rect -464 12 -444 14
rect -202 18 -182 20
rect -280 12 -260 14
rect -98 12 -78 14
rect -856 -37 -854 -17
rect -822 -38 -820 -18
rect -801 -38 -799 -18
rect -780 -38 -778 -18
rect -759 -38 -757 -18
rect -694 -30 -692 -10
rect -674 -30 -672 -10
rect -476 -34 -474 -14
rect -456 -34 -454 -14
rect -202 -2 -182 0
rect -292 -34 -290 -14
rect -272 -34 -270 -14
rect -110 -34 -108 -14
rect -90 -34 -88 -14
rect -553 -79 -551 -59
rect -532 -79 -530 -59
rect -511 -79 -509 -59
rect -369 -76 -367 -56
rect -348 -76 -346 -56
rect -327 -76 -325 -56
rect -809 -113 -789 -111
rect -731 -115 -729 -95
rect -710 -115 -708 -95
rect -689 -115 -687 -95
rect -668 -115 -666 -95
rect -638 -104 -636 -84
rect -617 -104 -615 -84
rect -596 -104 -594 -84
rect -809 -133 -789 -131
rect -462 -115 -460 -95
rect -441 -115 -439 -95
rect -420 -115 -418 -95
rect -399 -115 -397 -95
rect -596 -177 -576 -175
rect -596 -199 -576 -197
<< ndiffusion >>
rect -769 207 -759 208
rect -700 207 -690 208
rect -769 204 -759 205
rect -700 204 -690 205
rect -592 195 -582 196
rect -523 195 -513 196
rect -408 195 -398 196
rect -339 195 -329 196
rect -226 195 -216 196
rect -157 195 -147 196
rect -592 192 -582 193
rect -523 192 -513 193
rect -408 192 -398 193
rect -339 192 -329 193
rect -226 192 -216 193
rect -157 192 -147 193
rect -762 177 -752 178
rect -693 177 -683 178
rect -762 174 -752 175
rect -693 174 -683 175
rect -585 165 -575 166
rect -516 165 -506 166
rect -401 165 -391 166
rect -332 165 -322 166
rect -219 165 -209 166
rect -150 165 -140 166
rect -585 162 -575 163
rect -516 162 -506 163
rect -401 162 -391 163
rect -332 162 -322 163
rect -219 162 -209 163
rect -150 162 -140 163
rect -759 131 -758 141
rect -756 131 -755 141
rect -690 131 -689 141
rect -687 131 -686 141
rect -582 119 -581 129
rect -579 119 -578 129
rect -513 119 -512 129
rect -510 119 -509 129
rect -398 119 -397 129
rect -395 119 -394 129
rect -329 119 -328 129
rect -326 119 -325 129
rect -216 119 -215 129
rect -213 119 -212 129
rect -147 119 -146 129
rect -144 119 -143 129
rect -790 46 -789 56
rect -787 46 -786 56
rect -765 47 -764 87
rect -762 47 -761 87
rect -744 47 -743 87
rect -741 47 -740 87
rect -723 47 -722 87
rect -720 47 -719 87
rect -702 47 -701 87
rect -699 47 -698 87
rect -666 55 -665 75
rect -663 55 -662 75
rect -636 55 -635 75
rect -633 55 -632 75
rect -489 43 -488 63
rect -486 43 -485 63
rect -459 43 -458 63
rect -456 43 -455 63
rect -305 43 -304 63
rect -302 43 -301 63
rect -275 43 -274 63
rect -272 43 -271 63
rect -123 43 -122 63
rect -120 43 -119 63
rect -93 43 -92 63
rect -90 43 -89 63
rect -489 14 -479 15
rect -236 20 -216 21
rect -489 11 -479 12
rect -305 14 -295 15
rect -236 17 -216 18
rect -123 14 -113 15
rect -305 11 -295 12
rect -123 11 -113 12
rect -236 0 -216 1
rect -857 -62 -856 -52
rect -854 -62 -853 -52
rect -823 -93 -822 -53
rect -820 -93 -819 -53
rect -802 -93 -801 -53
rect -799 -93 -798 -53
rect -781 -93 -780 -53
rect -778 -93 -777 -53
rect -760 -93 -759 -53
rect -757 -93 -756 -53
rect -695 -64 -694 -44
rect -692 -64 -691 -44
rect -675 -64 -674 -44
rect -672 -64 -671 -44
rect -642 -48 -641 -8
rect -639 -48 -638 -8
rect -621 -48 -620 -8
rect -618 -48 -617 -8
rect -600 -48 -599 -8
rect -597 -48 -596 -8
rect -579 -48 -578 -8
rect -576 -48 -575 -8
rect -420 -30 -419 0
rect -417 -30 -416 0
rect -399 -30 -398 0
rect -396 -30 -395 0
rect -378 -30 -377 0
rect -375 -30 -374 0
rect -236 -3 -216 -2
rect -477 -68 -476 -48
rect -474 -68 -473 -48
rect -457 -68 -456 -48
rect -454 -68 -453 -48
rect -293 -68 -292 -48
rect -290 -68 -289 -48
rect -273 -68 -272 -48
rect -270 -68 -269 -48
rect -111 -68 -110 -48
rect -108 -68 -107 -48
rect -91 -68 -90 -48
rect -88 -68 -87 -48
rect -775 -111 -755 -110
rect -775 -114 -755 -113
rect -775 -131 -755 -130
rect -775 -134 -755 -133
rect -732 -170 -731 -130
rect -729 -170 -728 -130
rect -711 -170 -710 -130
rect -708 -170 -707 -130
rect -690 -170 -689 -130
rect -687 -170 -686 -130
rect -669 -170 -668 -130
rect -666 -170 -665 -130
rect -639 -149 -638 -119
rect -636 -149 -635 -119
rect -618 -149 -617 -119
rect -615 -149 -614 -119
rect -597 -149 -596 -119
rect -594 -149 -593 -119
rect -554 -124 -553 -94
rect -551 -124 -550 -94
rect -533 -124 -532 -94
rect -530 -124 -529 -94
rect -512 -124 -511 -94
rect -509 -124 -508 -94
rect -370 -121 -369 -91
rect -367 -121 -366 -91
rect -349 -121 -348 -91
rect -346 -121 -345 -91
rect -328 -121 -327 -91
rect -325 -121 -324 -91
rect -463 -170 -462 -130
rect -460 -170 -459 -130
rect -442 -170 -441 -130
rect -439 -170 -438 -130
rect -421 -170 -420 -130
rect -418 -170 -417 -130
rect -400 -170 -399 -130
rect -397 -170 -396 -130
rect -630 -175 -610 -174
rect -630 -178 -610 -177
rect -630 -197 -610 -196
rect -630 -200 -610 -199
<< pdiffusion >>
rect -744 207 -724 208
rect -672 207 -652 208
rect -744 204 -724 205
rect -672 204 -652 205
rect -567 195 -547 196
rect -495 195 -475 196
rect -383 195 -363 196
rect -311 195 -291 196
rect -201 195 -181 196
rect -129 195 -109 196
rect -567 192 -547 193
rect -495 192 -475 193
rect -383 192 -363 193
rect -311 192 -291 193
rect -201 192 -181 193
rect -129 192 -109 193
rect -737 177 -717 178
rect -665 177 -645 178
rect -737 174 -717 175
rect -665 174 -645 175
rect -560 165 -540 166
rect -488 165 -468 166
rect -376 165 -356 166
rect -304 165 -284 166
rect -194 165 -174 166
rect -122 165 -102 166
rect -560 162 -540 163
rect -488 162 -468 163
rect -376 162 -356 163
rect -304 162 -284 163
rect -194 162 -174 163
rect -122 162 -102 163
rect -733 131 -732 151
rect -730 131 -729 151
rect -661 131 -660 151
rect -658 131 -657 151
rect -556 119 -555 139
rect -553 119 -552 139
rect -484 119 -483 139
rect -481 119 -480 139
rect -372 119 -371 139
rect -369 119 -368 139
rect -300 119 -299 139
rect -297 119 -296 139
rect -190 119 -189 139
rect -187 119 -186 139
rect -118 119 -117 139
rect -115 119 -114 139
rect -666 89 -665 109
rect -663 89 -662 109
rect -636 89 -635 109
rect -633 89 -632 109
rect -489 77 -488 97
rect -486 77 -485 97
rect -459 77 -458 97
rect -456 77 -455 97
rect -305 77 -304 97
rect -302 77 -301 97
rect -275 77 -274 97
rect -272 77 -271 97
rect -123 77 -122 97
rect -120 77 -119 97
rect -93 77 -92 97
rect -90 77 -89 97
rect -790 12 -789 32
rect -787 12 -786 32
rect -765 12 -764 32
rect -762 12 -761 32
rect -744 12 -743 32
rect -741 12 -740 32
rect -723 12 -722 32
rect -720 12 -719 32
rect -702 12 -701 32
rect -699 12 -698 32
rect -642 7 -641 27
rect -639 7 -638 27
rect -621 7 -620 27
rect -618 7 -617 27
rect -600 7 -599 27
rect -597 7 -596 27
rect -579 7 -578 27
rect -576 7 -575 27
rect -420 15 -419 35
rect -417 15 -416 35
rect -399 15 -398 35
rect -396 15 -395 35
rect -378 15 -377 35
rect -375 15 -374 35
rect -202 20 -182 21
rect -464 14 -444 15
rect -464 11 -444 12
rect -280 14 -260 15
rect -202 17 -182 18
rect -98 14 -78 15
rect -280 11 -260 12
rect -98 11 -78 12
rect -202 0 -182 1
rect -857 -37 -856 -17
rect -854 -37 -853 -17
rect -823 -38 -822 -18
rect -820 -38 -819 -18
rect -802 -38 -801 -18
rect -799 -38 -798 -18
rect -781 -38 -780 -18
rect -778 -38 -777 -18
rect -760 -38 -759 -18
rect -757 -38 -756 -18
rect -695 -30 -694 -10
rect -692 -30 -691 -10
rect -675 -30 -674 -10
rect -672 -30 -671 -10
rect -477 -34 -476 -14
rect -474 -34 -473 -14
rect -457 -34 -456 -14
rect -454 -34 -453 -14
rect -202 -3 -182 -2
rect -293 -34 -292 -14
rect -290 -34 -289 -14
rect -273 -34 -272 -14
rect -270 -34 -269 -14
rect -111 -34 -110 -14
rect -108 -34 -107 -14
rect -91 -34 -90 -14
rect -88 -34 -87 -14
rect -554 -79 -553 -59
rect -551 -79 -550 -59
rect -533 -79 -532 -59
rect -530 -79 -529 -59
rect -512 -79 -511 -59
rect -509 -79 -508 -59
rect -370 -76 -369 -56
rect -367 -76 -366 -56
rect -349 -76 -348 -56
rect -346 -76 -345 -56
rect -328 -76 -327 -56
rect -325 -76 -324 -56
rect -809 -111 -789 -110
rect -809 -114 -789 -113
rect -732 -115 -731 -95
rect -729 -115 -728 -95
rect -711 -115 -710 -95
rect -708 -115 -707 -95
rect -690 -115 -689 -95
rect -687 -115 -686 -95
rect -669 -115 -668 -95
rect -666 -115 -665 -95
rect -639 -104 -638 -84
rect -636 -104 -635 -84
rect -618 -104 -617 -84
rect -615 -104 -614 -84
rect -597 -104 -596 -84
rect -594 -104 -593 -84
rect -809 -131 -789 -130
rect -809 -134 -789 -133
rect -463 -115 -462 -95
rect -460 -115 -459 -95
rect -442 -115 -441 -95
rect -439 -115 -438 -95
rect -421 -115 -420 -95
rect -418 -115 -417 -95
rect -400 -115 -399 -95
rect -397 -115 -396 -95
rect -596 -175 -576 -174
rect -596 -178 -576 -177
rect -596 -197 -576 -196
rect -596 -200 -576 -199
<< ndcontact >>
rect -769 208 -759 212
rect -700 208 -690 212
rect -769 200 -759 204
rect -700 200 -690 204
rect -592 196 -582 200
rect -523 196 -513 200
rect -408 196 -398 200
rect -339 196 -329 200
rect -226 196 -216 200
rect -157 196 -147 200
rect -592 188 -582 192
rect -523 188 -513 192
rect -408 188 -398 192
rect -339 188 -329 192
rect -226 188 -216 192
rect -157 188 -147 192
rect -762 178 -752 182
rect -693 178 -683 182
rect -762 170 -752 174
rect -693 170 -683 174
rect -585 166 -575 170
rect -516 166 -506 170
rect -401 166 -391 170
rect -332 166 -322 170
rect -219 166 -209 170
rect -150 166 -140 170
rect -585 158 -575 162
rect -516 158 -506 162
rect -401 158 -391 162
rect -332 158 -322 162
rect -219 158 -209 162
rect -150 158 -140 162
rect -763 131 -759 141
rect -755 131 -751 141
rect -694 131 -690 141
rect -686 131 -682 141
rect -586 119 -582 129
rect -578 119 -574 129
rect -517 119 -513 129
rect -509 119 -505 129
rect -402 119 -398 129
rect -394 119 -390 129
rect -333 119 -329 129
rect -325 119 -321 129
rect -220 119 -216 129
rect -212 119 -208 129
rect -151 119 -147 129
rect -143 119 -139 129
rect -794 46 -790 56
rect -786 46 -782 56
rect -769 47 -765 87
rect -761 47 -757 87
rect -748 47 -744 87
rect -740 47 -736 87
rect -727 47 -723 87
rect -719 47 -715 87
rect -706 47 -702 87
rect -698 47 -694 87
rect -670 55 -666 75
rect -662 55 -658 75
rect -640 55 -636 75
rect -632 55 -628 75
rect -493 43 -489 63
rect -485 43 -481 63
rect -463 43 -459 63
rect -455 43 -451 63
rect -309 43 -305 63
rect -301 43 -297 63
rect -279 43 -275 63
rect -271 43 -267 63
rect -127 43 -123 63
rect -119 43 -115 63
rect -97 43 -93 63
rect -89 43 -85 63
rect -489 15 -479 19
rect -236 21 -216 25
rect -305 15 -295 19
rect -489 7 -479 11
rect -236 13 -216 17
rect -123 15 -113 19
rect -305 7 -295 11
rect -123 7 -113 11
rect -236 1 -216 5
rect -861 -62 -857 -52
rect -853 -62 -849 -52
rect -827 -93 -823 -53
rect -819 -93 -815 -53
rect -806 -93 -802 -53
rect -798 -93 -794 -53
rect -785 -93 -781 -53
rect -777 -93 -773 -53
rect -764 -93 -760 -53
rect -756 -93 -752 -53
rect -699 -64 -695 -44
rect -691 -64 -687 -44
rect -679 -64 -675 -44
rect -671 -64 -667 -44
rect -646 -48 -642 -8
rect -638 -48 -634 -8
rect -625 -48 -621 -8
rect -617 -48 -613 -8
rect -604 -48 -600 -8
rect -596 -48 -592 -8
rect -583 -48 -579 -8
rect -575 -48 -571 -8
rect -424 -30 -420 0
rect -416 -30 -412 0
rect -403 -30 -399 0
rect -395 -30 -391 0
rect -382 -30 -378 0
rect -374 -30 -370 0
rect -236 -7 -216 -3
rect -481 -68 -477 -48
rect -473 -68 -469 -48
rect -461 -68 -457 -48
rect -453 -68 -449 -48
rect -297 -68 -293 -48
rect -289 -68 -285 -48
rect -277 -68 -273 -48
rect -269 -68 -265 -48
rect -115 -68 -111 -48
rect -107 -68 -103 -48
rect -95 -68 -91 -48
rect -87 -68 -83 -48
rect -775 -110 -755 -106
rect -775 -118 -755 -114
rect -775 -130 -755 -126
rect -775 -138 -755 -134
rect -736 -170 -732 -130
rect -728 -170 -724 -130
rect -715 -170 -711 -130
rect -707 -170 -703 -130
rect -694 -170 -690 -130
rect -686 -170 -682 -130
rect -673 -170 -669 -130
rect -665 -170 -661 -130
rect -643 -149 -639 -119
rect -635 -149 -631 -119
rect -622 -149 -618 -119
rect -614 -149 -610 -119
rect -601 -149 -597 -119
rect -593 -149 -589 -119
rect -558 -124 -554 -94
rect -550 -124 -546 -94
rect -537 -124 -533 -94
rect -529 -124 -525 -94
rect -516 -124 -512 -94
rect -508 -124 -504 -94
rect -374 -121 -370 -91
rect -366 -121 -362 -91
rect -353 -121 -349 -91
rect -345 -121 -341 -91
rect -332 -121 -328 -91
rect -324 -121 -320 -91
rect -467 -170 -463 -130
rect -459 -170 -455 -130
rect -446 -170 -442 -130
rect -438 -170 -434 -130
rect -425 -170 -421 -130
rect -417 -170 -413 -130
rect -404 -170 -400 -130
rect -396 -170 -392 -130
rect -630 -174 -610 -170
rect -630 -182 -610 -178
rect -630 -196 -610 -192
rect -630 -204 -610 -200
<< pdcontact >>
rect -744 208 -724 212
rect -672 208 -652 212
rect -744 200 -724 204
rect -672 200 -652 204
rect -567 196 -547 200
rect -495 196 -475 200
rect -383 196 -363 200
rect -311 196 -291 200
rect -201 196 -181 200
rect -129 196 -109 200
rect -567 188 -547 192
rect -495 188 -475 192
rect -383 188 -363 192
rect -311 188 -291 192
rect -201 188 -181 192
rect -129 188 -109 192
rect -737 178 -717 182
rect -665 178 -645 182
rect -737 170 -717 174
rect -665 170 -645 174
rect -560 166 -540 170
rect -488 166 -468 170
rect -376 166 -356 170
rect -304 166 -284 170
rect -194 166 -174 170
rect -122 166 -102 170
rect -560 158 -540 162
rect -488 158 -468 162
rect -376 158 -356 162
rect -304 158 -284 162
rect -194 158 -174 162
rect -122 158 -102 162
rect -737 131 -733 151
rect -729 131 -725 151
rect -665 131 -661 151
rect -657 131 -653 151
rect -560 119 -556 139
rect -552 119 -548 139
rect -488 119 -484 139
rect -480 119 -476 139
rect -376 119 -372 139
rect -368 119 -364 139
rect -304 119 -300 139
rect -296 119 -292 139
rect -194 119 -190 139
rect -186 119 -182 139
rect -122 119 -118 139
rect -114 119 -110 139
rect -670 89 -666 109
rect -662 89 -658 109
rect -640 89 -636 109
rect -632 89 -628 109
rect -493 77 -489 97
rect -485 77 -481 97
rect -463 77 -459 97
rect -455 77 -451 97
rect -309 77 -305 97
rect -301 77 -297 97
rect -279 77 -275 97
rect -271 77 -267 97
rect -127 77 -123 97
rect -119 77 -115 97
rect -97 77 -93 97
rect -89 77 -85 97
rect -794 12 -790 32
rect -786 12 -782 32
rect -769 12 -765 32
rect -761 12 -757 32
rect -748 12 -744 32
rect -740 12 -736 32
rect -727 12 -723 32
rect -719 12 -715 32
rect -706 12 -702 32
rect -698 12 -694 32
rect -646 7 -642 27
rect -638 7 -634 27
rect -625 7 -621 27
rect -617 7 -613 27
rect -604 7 -600 27
rect -596 7 -592 27
rect -583 7 -579 27
rect -575 7 -571 27
rect -464 15 -444 19
rect -424 15 -420 35
rect -416 15 -412 35
rect -403 15 -399 35
rect -395 15 -391 35
rect -382 15 -378 35
rect -374 15 -370 35
rect -202 21 -182 25
rect -464 7 -444 11
rect -280 15 -260 19
rect -202 13 -182 17
rect -98 15 -78 19
rect -280 7 -260 11
rect -98 7 -78 11
rect -202 1 -182 5
rect -861 -37 -857 -17
rect -853 -37 -849 -17
rect -827 -38 -823 -18
rect -819 -38 -815 -18
rect -806 -38 -802 -18
rect -798 -38 -794 -18
rect -785 -38 -781 -18
rect -777 -38 -773 -18
rect -764 -38 -760 -18
rect -756 -38 -752 -18
rect -699 -30 -695 -10
rect -691 -30 -687 -10
rect -679 -30 -675 -10
rect -671 -30 -667 -10
rect -481 -34 -477 -14
rect -473 -34 -469 -14
rect -461 -34 -457 -14
rect -453 -34 -449 -14
rect -202 -7 -182 -3
rect -297 -34 -293 -14
rect -289 -34 -285 -14
rect -277 -34 -273 -14
rect -269 -34 -265 -14
rect -115 -34 -111 -14
rect -107 -34 -103 -14
rect -95 -34 -91 -14
rect -87 -34 -83 -14
rect -558 -79 -554 -59
rect -550 -79 -546 -59
rect -537 -79 -533 -59
rect -529 -79 -525 -59
rect -516 -79 -512 -59
rect -508 -79 -504 -59
rect -374 -76 -370 -56
rect -366 -76 -362 -56
rect -353 -76 -349 -56
rect -345 -76 -341 -56
rect -332 -76 -328 -56
rect -324 -76 -320 -56
rect -809 -110 -789 -106
rect -809 -118 -789 -114
rect -736 -115 -732 -95
rect -728 -115 -724 -95
rect -715 -115 -711 -95
rect -707 -115 -703 -95
rect -694 -115 -690 -95
rect -686 -115 -682 -95
rect -673 -115 -669 -95
rect -665 -115 -661 -95
rect -643 -104 -639 -84
rect -635 -104 -631 -84
rect -622 -104 -618 -84
rect -614 -104 -610 -84
rect -601 -104 -597 -84
rect -593 -104 -589 -84
rect -809 -130 -789 -126
rect -809 -138 -789 -134
rect -467 -115 -463 -95
rect -459 -115 -455 -95
rect -446 -115 -442 -95
rect -438 -115 -434 -95
rect -425 -115 -421 -95
rect -417 -115 -413 -95
rect -404 -115 -400 -95
rect -396 -115 -392 -95
rect -596 -174 -576 -170
rect -596 -182 -576 -178
rect -596 -196 -576 -192
rect -596 -204 -576 -200
<< polysilicon >>
rect -772 205 -769 207
rect -759 205 -744 207
rect -724 205 -721 207
rect -703 205 -700 207
rect -690 205 -672 207
rect -652 205 -649 207
rect -595 193 -592 195
rect -582 193 -567 195
rect -547 193 -544 195
rect -526 193 -523 195
rect -513 193 -495 195
rect -475 193 -472 195
rect -411 193 -408 195
rect -398 193 -383 195
rect -363 193 -360 195
rect -342 193 -339 195
rect -329 193 -311 195
rect -291 193 -288 195
rect -229 193 -226 195
rect -216 193 -201 195
rect -181 193 -178 195
rect -160 193 -157 195
rect -147 193 -129 195
rect -109 193 -106 195
rect -765 175 -762 177
rect -752 175 -737 177
rect -717 175 -714 177
rect -696 175 -693 177
rect -683 175 -665 177
rect -645 175 -642 177
rect -588 163 -585 165
rect -575 163 -560 165
rect -540 163 -537 165
rect -519 163 -516 165
rect -506 163 -488 165
rect -468 163 -465 165
rect -404 163 -401 165
rect -391 163 -376 165
rect -356 163 -353 165
rect -335 163 -332 165
rect -322 163 -304 165
rect -284 163 -281 165
rect -222 163 -219 165
rect -209 163 -194 165
rect -174 163 -171 165
rect -153 163 -150 165
rect -140 163 -122 165
rect -102 163 -99 165
rect -732 151 -730 163
rect -660 151 -658 163
rect -758 141 -756 148
rect -689 141 -687 148
rect -555 139 -553 151
rect -483 139 -481 151
rect -371 139 -369 151
rect -299 139 -297 151
rect -189 139 -187 151
rect -117 139 -115 151
rect -758 128 -756 131
rect -732 128 -730 131
rect -689 128 -687 131
rect -660 128 -658 131
rect -581 129 -579 136
rect -512 129 -510 136
rect -397 129 -395 136
rect -328 129 -326 136
rect -215 129 -213 136
rect -146 129 -144 136
rect -581 116 -579 119
rect -555 116 -553 119
rect -512 116 -510 119
rect -483 116 -481 119
rect -397 116 -395 119
rect -371 116 -369 119
rect -328 116 -326 119
rect -299 116 -297 119
rect -215 116 -213 119
rect -189 116 -187 119
rect -146 116 -144 119
rect -117 116 -115 119
rect -665 109 -663 112
rect -635 109 -633 112
rect -764 87 -762 91
rect -743 87 -741 91
rect -722 87 -720 91
rect -701 87 -699 91
rect -488 97 -486 100
rect -458 97 -456 100
rect -304 97 -302 100
rect -274 97 -272 100
rect -122 97 -120 100
rect -92 97 -90 100
rect -789 56 -787 59
rect -665 75 -663 89
rect -635 75 -633 89
rect -488 63 -486 77
rect -458 63 -456 77
rect -304 63 -302 77
rect -274 63 -272 77
rect -122 63 -120 77
rect -92 63 -90 77
rect -665 51 -663 55
rect -635 51 -633 55
rect -789 32 -787 46
rect -764 32 -762 47
rect -743 32 -741 47
rect -722 32 -720 47
rect -701 32 -699 47
rect -488 39 -486 43
rect -458 39 -456 43
rect -304 39 -302 43
rect -274 39 -272 43
rect -122 39 -120 43
rect -92 39 -90 43
rect -419 35 -417 38
rect -398 35 -396 38
rect -377 35 -375 38
rect -641 27 -639 30
rect -620 27 -618 30
rect -599 27 -597 30
rect -578 27 -576 30
rect -789 9 -787 12
rect -764 9 -762 12
rect -743 9 -741 12
rect -722 9 -720 12
rect -701 9 -699 12
rect -492 12 -489 14
rect -479 12 -464 14
rect -444 12 -441 14
rect -694 -10 -692 -7
rect -674 -10 -672 -7
rect -641 -8 -639 7
rect -620 -8 -618 7
rect -599 -8 -597 7
rect -578 -8 -576 7
rect -419 0 -417 15
rect -398 0 -396 15
rect -377 0 -375 15
rect -240 18 -236 20
rect -216 18 -202 20
rect -182 18 -179 20
rect -308 12 -305 14
rect -295 12 -280 14
rect -260 12 -257 14
rect -126 12 -123 14
rect -113 12 -98 14
rect -78 12 -75 14
rect -856 -17 -854 -14
rect -822 -18 -820 -15
rect -801 -18 -799 -15
rect -780 -18 -778 -15
rect -759 -18 -757 -15
rect -856 -52 -854 -37
rect -822 -53 -820 -38
rect -801 -53 -799 -38
rect -780 -53 -778 -38
rect -759 -53 -757 -38
rect -694 -44 -692 -30
rect -674 -44 -672 -30
rect -856 -65 -854 -62
rect -476 -14 -474 -11
rect -456 -14 -454 -11
rect -240 -2 -236 0
rect -216 -2 -202 0
rect -182 -2 -179 0
rect -292 -14 -290 -11
rect -272 -14 -270 -11
rect -110 -14 -108 -11
rect -90 -14 -88 -11
rect -419 -34 -417 -30
rect -398 -34 -396 -30
rect -377 -34 -375 -30
rect -476 -48 -474 -34
rect -456 -48 -454 -34
rect -292 -48 -290 -34
rect -272 -48 -270 -34
rect -110 -48 -108 -34
rect -90 -48 -88 -34
rect -641 -52 -639 -48
rect -620 -52 -618 -48
rect -599 -52 -597 -48
rect -578 -52 -576 -48
rect -553 -59 -551 -56
rect -532 -59 -530 -56
rect -511 -59 -509 -56
rect -694 -68 -692 -64
rect -674 -68 -672 -64
rect -369 -56 -367 -53
rect -348 -56 -346 -53
rect -327 -56 -325 -53
rect -476 -72 -474 -68
rect -456 -71 -454 -68
rect -292 -72 -290 -68
rect -272 -72 -270 -68
rect -110 -72 -108 -68
rect -90 -72 -88 -68
rect -638 -84 -636 -81
rect -617 -84 -615 -81
rect -596 -84 -594 -81
rect -822 -97 -820 -93
rect -801 -97 -799 -93
rect -780 -97 -778 -93
rect -759 -97 -757 -93
rect -731 -95 -729 -92
rect -710 -95 -708 -92
rect -689 -95 -687 -92
rect -668 -95 -666 -92
rect -812 -113 -809 -111
rect -789 -113 -775 -111
rect -755 -113 -751 -111
rect -553 -94 -551 -79
rect -532 -94 -530 -79
rect -511 -94 -509 -79
rect -369 -91 -367 -76
rect -348 -91 -346 -76
rect -327 -91 -325 -76
rect -731 -130 -729 -115
rect -710 -130 -708 -115
rect -689 -130 -687 -115
rect -668 -130 -666 -115
rect -638 -119 -636 -104
rect -617 -119 -615 -104
rect -596 -119 -594 -104
rect -812 -133 -809 -131
rect -789 -133 -775 -131
rect -755 -133 -751 -131
rect -462 -95 -460 -92
rect -441 -95 -439 -92
rect -420 -95 -418 -92
rect -399 -95 -397 -92
rect -553 -128 -551 -124
rect -532 -128 -530 -124
rect -511 -128 -509 -124
rect -462 -130 -460 -115
rect -441 -130 -439 -115
rect -420 -130 -418 -115
rect -399 -130 -397 -115
rect -369 -125 -367 -121
rect -348 -125 -346 -121
rect -327 -125 -325 -121
rect -638 -153 -636 -149
rect -617 -153 -615 -149
rect -596 -153 -594 -149
rect -731 -174 -729 -170
rect -710 -174 -708 -170
rect -689 -174 -687 -170
rect -668 -174 -666 -170
rect -462 -174 -460 -170
rect -441 -174 -439 -170
rect -420 -174 -418 -170
rect -399 -174 -397 -170
rect -634 -177 -630 -175
rect -610 -177 -596 -175
rect -576 -177 -573 -175
rect -634 -199 -630 -197
rect -610 -199 -596 -197
rect -576 -199 -573 -197
<< polycontact >>
rect -756 207 -752 211
rect -687 207 -683 211
rect -579 195 -575 199
rect -510 195 -506 199
rect -395 195 -391 199
rect -326 195 -322 199
rect -213 195 -209 199
rect -144 195 -140 199
rect -749 177 -745 181
rect -677 177 -673 181
rect -572 165 -568 169
rect -500 165 -496 169
rect -388 165 -384 169
rect -316 165 -312 169
rect -206 165 -202 169
rect -134 165 -130 169
rect -730 159 -726 163
rect -658 159 -654 163
rect -762 144 -758 148
rect -693 144 -689 148
rect -553 147 -549 151
rect -481 147 -477 151
rect -369 147 -365 151
rect -297 147 -293 151
rect -187 147 -183 151
rect -115 147 -111 151
rect -585 132 -581 136
rect -516 132 -512 136
rect -401 132 -397 136
rect -332 132 -328 136
rect -219 132 -215 136
rect -150 132 -146 136
rect -669 78 -665 82
rect -633 78 -629 82
rect -492 66 -488 70
rect -456 66 -452 70
rect -308 66 -304 70
rect -272 66 -268 70
rect -126 66 -122 70
rect -90 66 -86 70
rect -787 39 -783 43
rect -762 39 -758 43
rect -741 39 -737 43
rect -720 39 -716 43
rect -699 39 -695 43
rect -476 14 -472 18
rect -213 20 -209 24
rect -639 -4 -635 0
rect -618 -4 -614 0
rect -597 -4 -593 0
rect -417 4 -413 8
rect -396 4 -392 8
rect -292 14 -288 18
rect -110 14 -106 18
rect -375 4 -371 8
rect -576 -4 -572 0
rect -854 -49 -850 -45
rect -820 -49 -816 -45
rect -799 -49 -795 -45
rect -778 -49 -774 -45
rect -698 -41 -694 -37
rect -672 -41 -668 -37
rect -757 -49 -753 -45
rect -213 -6 -209 -2
rect -480 -45 -476 -41
rect -454 -45 -450 -41
rect -296 -45 -292 -41
rect -270 -45 -266 -41
rect -114 -45 -110 -41
rect -88 -45 -84 -41
rect -782 -111 -778 -107
rect -551 -90 -547 -86
rect -530 -90 -526 -86
rect -509 -90 -505 -86
rect -367 -87 -363 -83
rect -346 -87 -342 -83
rect -325 -87 -321 -83
rect -729 -126 -725 -122
rect -708 -126 -704 -122
rect -687 -126 -683 -122
rect -636 -115 -632 -111
rect -615 -115 -611 -111
rect -594 -115 -590 -111
rect -666 -126 -662 -122
rect -782 -137 -778 -133
rect -460 -126 -456 -122
rect -439 -126 -435 -122
rect -418 -126 -414 -122
rect -397 -126 -393 -122
rect -607 -175 -603 -171
rect -607 -203 -603 -199
<< metal1 >>
rect -756 221 -708 225
rect -773 208 -769 212
rect -756 211 -752 221
rect -720 212 -716 218
rect -724 208 -716 212
rect -759 200 -744 204
rect -756 197 -752 200
rect -770 194 -752 197
rect -720 198 -716 208
rect -770 182 -766 194
rect -770 178 -762 182
rect -749 181 -745 185
rect -712 182 -708 221
rect -687 221 -636 225
rect -687 211 -683 221
rect -648 212 -644 218
rect -652 208 -644 212
rect -690 200 -672 204
rect -687 197 -683 200
rect -770 148 -766 178
rect -717 178 -708 182
rect -752 170 -737 174
rect -749 163 -745 170
rect -712 163 -708 178
rect -754 160 -733 163
rect -754 158 -751 160
rect -770 144 -762 148
rect -755 141 -751 158
rect -737 151 -733 160
rect -726 159 -713 163
rect -763 127 -759 131
rect -729 127 -725 131
rect -763 123 -750 127
rect -745 123 -719 127
rect -713 119 -708 158
rect -701 194 -683 197
rect -648 198 -644 208
rect -640 207 -636 221
rect -579 209 -531 213
rect -701 182 -697 194
rect -652 193 -648 196
rect -701 178 -693 182
rect -677 181 -673 185
rect -640 182 -636 202
rect -596 196 -592 200
rect -579 199 -575 209
rect -543 200 -539 206
rect -547 196 -539 200
rect -582 188 -567 192
rect -579 185 -575 188
rect -701 148 -697 178
rect -645 178 -636 182
rect -593 182 -575 185
rect -543 186 -539 196
rect -683 170 -665 174
rect -677 163 -673 170
rect -640 163 -636 178
rect -682 160 -661 163
rect -701 144 -693 148
rect -686 141 -682 158
rect -665 151 -661 160
rect -654 159 -636 163
rect -593 170 -589 182
rect -593 166 -585 170
rect -572 169 -568 173
rect -535 170 -531 209
rect -510 209 -459 213
rect -510 199 -506 209
rect -471 200 -467 206
rect -475 196 -467 200
rect -513 188 -495 192
rect -510 185 -506 188
rect -593 136 -589 166
rect -540 166 -531 170
rect -575 158 -560 162
rect -572 151 -568 158
rect -535 151 -531 166
rect -577 148 -556 151
rect -577 146 -574 148
rect -593 132 -585 136
rect -694 127 -690 131
rect -657 127 -653 131
rect -578 129 -574 146
rect -694 123 -678 127
rect -673 123 -647 127
rect -560 139 -556 148
rect -549 147 -536 151
rect -713 116 -685 119
rect -780 65 -777 92
rect -761 88 -744 91
rect -761 87 -757 88
rect -786 61 -777 65
rect -786 56 -783 61
rect -748 87 -744 88
rect -740 88 -723 91
rect -740 87 -736 88
rect -727 87 -723 88
rect -719 88 -702 91
rect -719 87 -715 88
rect -706 87 -702 88
rect -698 87 -694 92
rect -794 43 -790 46
rect -797 40 -790 43
rect -794 32 -790 40
rect -783 39 -779 43
rect -769 43 -765 47
rect -688 44 -685 116
rect -676 113 -652 117
rect -646 113 -622 117
rect -586 115 -582 119
rect -552 115 -548 119
rect -670 109 -666 113
rect -632 109 -628 113
rect -586 111 -573 115
rect -662 82 -658 89
rect -568 111 -542 115
rect -640 82 -636 89
rect -673 78 -669 82
rect -662 78 -653 82
rect -648 78 -636 82
rect -629 78 -625 82
rect -640 75 -636 78
rect -670 50 -666 55
rect -669 46 -666 50
rect -573 61 -568 110
rect -662 50 -658 55
rect -632 50 -628 55
rect -662 46 -628 50
rect -774 39 -765 43
rect -690 41 -685 44
rect -769 32 -765 39
rect -748 32 -744 39
rect -727 32 -723 39
rect -706 32 -702 39
rect -536 35 -531 146
rect -524 182 -506 185
rect -471 186 -467 196
rect -463 195 -459 209
rect -395 209 -347 213
rect -412 196 -408 200
rect -395 199 -391 209
rect -359 200 -355 206
rect -363 196 -355 200
rect -524 170 -520 182
rect -475 181 -471 184
rect -524 166 -516 170
rect -500 169 -496 173
rect -463 170 -459 190
rect -398 188 -383 192
rect -395 185 -391 188
rect -409 182 -391 185
rect -359 186 -355 196
rect -524 136 -520 166
rect -468 166 -459 170
rect -506 158 -488 162
rect -500 151 -496 158
rect -463 151 -459 166
rect -505 148 -484 151
rect -524 132 -516 136
rect -509 129 -505 146
rect -488 139 -484 148
rect -477 147 -459 151
rect -409 170 -405 182
rect -409 166 -401 170
rect -388 169 -384 173
rect -351 170 -347 209
rect -326 209 -275 213
rect -326 199 -322 209
rect -287 200 -283 206
rect -291 196 -283 200
rect -329 188 -311 192
rect -326 185 -322 188
rect -409 136 -405 166
rect -356 166 -347 170
rect -391 158 -376 162
rect -388 151 -384 158
rect -351 151 -347 166
rect -393 148 -372 151
rect -393 146 -390 148
rect -409 132 -401 136
rect -394 129 -390 146
rect -517 115 -513 119
rect -480 115 -476 119
rect -376 139 -372 148
rect -365 147 -352 151
rect -402 115 -398 119
rect -368 115 -364 119
rect -517 111 -501 115
rect -496 111 -470 115
rect -402 111 -389 115
rect -384 111 -358 115
rect -508 101 -475 105
rect -469 101 -445 105
rect -652 34 -565 35
rect -786 8 -782 12
rect -761 8 -757 12
rect -740 8 -736 12
rect -719 8 -715 12
rect -698 8 -694 12
rect -676 31 -550 34
rect -536 32 -511 35
rect -676 8 -673 31
rect -638 27 -634 31
rect -617 27 -613 31
rect -596 27 -592 31
rect -575 27 -571 31
rect -800 5 -673 8
rect -800 4 -688 5
rect -867 -10 -843 -9
rect -800 -10 -797 4
rect -676 -2 -673 5
rect -646 0 -642 7
rect -625 0 -621 7
rect -604 0 -600 7
rect -583 0 -579 7
rect -712 -5 -661 -2
rect -572 -4 -562 -1
rect -867 -13 -746 -10
rect -853 -17 -849 -13
rect -836 -14 -746 -13
rect -861 -45 -857 -37
rect -864 -49 -857 -45
rect -850 -49 -846 -45
rect -861 -52 -857 -49
rect -853 -63 -849 -62
rect -836 -100 -833 -14
rect -819 -18 -815 -14
rect -798 -18 -794 -14
rect -777 -18 -773 -14
rect -756 -18 -752 -14
rect -827 -45 -823 -38
rect -806 -45 -802 -38
rect -785 -45 -781 -38
rect -764 -45 -760 -38
rect -753 -49 -744 -46
rect -827 -53 -823 -50
rect -747 -53 -744 -49
rect -819 -94 -815 -93
rect -806 -94 -802 -93
rect -819 -97 -802 -94
rect -798 -94 -794 -93
rect -785 -94 -781 -93
rect -798 -97 -781 -94
rect -777 -94 -773 -93
rect -764 -94 -760 -93
rect -777 -97 -760 -94
rect -756 -94 -752 -93
rect -712 -76 -709 -5
rect -705 -6 -661 -5
rect -699 -10 -695 -6
rect -671 -10 -667 -6
rect -646 -8 -642 -5
rect -691 -36 -687 -30
rect -650 -14 -649 -11
rect -700 -41 -698 -37
rect -691 -40 -684 -36
rect -691 -44 -687 -40
rect -679 -40 -675 -30
rect -699 -69 -695 -64
rect -679 -69 -675 -64
rect -699 -73 -675 -69
rect -652 -55 -649 -14
rect -638 -49 -634 -48
rect -625 -49 -621 -48
rect -638 -52 -621 -49
rect -617 -49 -613 -48
rect -604 -49 -600 -48
rect -617 -52 -600 -49
rect -596 -49 -592 -48
rect -583 -49 -579 -48
rect -596 -52 -579 -49
rect -575 -49 -571 -48
rect -553 -51 -550 31
rect -514 -41 -511 32
rect -508 -5 -504 101
rect -493 97 -489 101
rect -455 97 -451 101
rect -485 70 -481 77
rect -463 70 -459 77
rect -496 66 -492 70
rect -485 66 -476 70
rect -471 66 -459 70
rect -452 66 -448 70
rect -493 40 -489 43
rect -492 35 -489 40
rect -485 37 -481 43
rect -476 45 -471 65
rect -463 63 -459 66
rect -389 61 -384 110
rect -455 37 -451 43
rect -430 39 -368 43
rect -497 20 -493 35
rect -485 34 -451 37
rect -416 35 -412 39
rect -395 35 -391 39
rect -374 35 -370 39
rect -493 15 -489 19
rect -476 18 -472 26
rect -440 19 -436 25
rect -444 15 -436 19
rect -479 7 -464 11
rect -476 2 -472 7
rect -503 -10 -448 -6
rect -440 -6 -436 15
rect -424 8 -420 15
rect -403 8 -399 15
rect -382 8 -378 15
rect -443 -10 -436 -6
rect -424 0 -420 3
rect -481 -14 -477 -10
rect -453 -14 -449 -10
rect -514 -43 -480 -41
rect -542 -45 -480 -43
rect -473 -44 -469 -34
rect -416 -31 -412 -30
rect -403 -31 -399 -30
rect -416 -34 -399 -31
rect -395 -31 -391 -30
rect -382 -31 -378 -30
rect -461 -41 -457 -34
rect -395 -35 -378 -31
rect -374 -31 -370 -30
rect -352 -38 -347 146
rect -340 182 -322 185
rect -287 186 -283 196
rect -279 195 -275 209
rect -213 209 -165 213
rect -230 196 -226 200
rect -213 199 -209 209
rect -177 200 -173 206
rect -181 196 -173 200
rect -340 170 -336 182
rect -291 181 -287 184
rect -340 166 -332 170
rect -316 169 -312 173
rect -279 170 -275 190
rect -216 188 -201 192
rect -213 185 -209 188
rect -227 182 -209 185
rect -177 186 -173 196
rect -340 136 -336 166
rect -284 166 -275 170
rect -322 158 -304 162
rect -316 151 -312 158
rect -279 151 -275 166
rect -321 148 -300 151
rect -340 132 -332 136
rect -325 129 -321 146
rect -304 139 -300 148
rect -293 147 -275 151
rect -227 170 -223 182
rect -227 166 -219 170
rect -206 169 -202 173
rect -169 170 -165 209
rect -144 209 -93 213
rect -144 199 -140 209
rect -105 200 -101 206
rect -109 196 -101 200
rect -147 188 -129 192
rect -144 185 -140 188
rect -227 136 -223 166
rect -174 166 -165 170
rect -209 158 -194 162
rect -206 151 -202 158
rect -169 151 -165 166
rect -211 148 -190 151
rect -211 146 -208 148
rect -227 132 -219 136
rect -212 129 -208 146
rect -333 115 -329 119
rect -296 115 -292 119
rect -194 139 -190 148
rect -183 147 -170 151
rect -158 182 -140 185
rect -105 186 -101 196
rect -97 195 -93 209
rect -158 170 -154 182
rect -109 181 -105 184
rect -158 166 -150 170
rect -134 169 -130 173
rect -97 170 -93 190
rect -220 115 -216 119
rect -186 115 -182 119
rect -333 111 -317 115
rect -312 111 -286 115
rect -220 111 -207 115
rect -202 111 -176 115
rect -324 101 -291 105
rect -285 101 -261 105
rect -324 45 -320 101
rect -309 97 -305 101
rect -271 97 -267 101
rect -301 70 -297 77
rect -279 70 -275 77
rect -312 66 -308 70
rect -301 66 -292 70
rect -287 66 -275 70
rect -268 66 -264 70
rect -332 3 -329 31
rect -324 -6 -320 40
rect -309 38 -305 43
rect -308 34 -305 38
rect -301 37 -297 43
rect -292 45 -287 65
rect -279 63 -275 66
rect -207 61 -202 110
rect -271 37 -267 43
rect -301 34 -267 37
rect -313 20 -309 33
rect -309 15 -305 19
rect -292 18 -288 26
rect -256 19 -252 25
rect -213 24 -209 26
rect -178 25 -174 31
rect -182 21 -174 25
rect -260 15 -252 19
rect -295 7 -293 11
rect -288 7 -280 11
rect -256 -6 -252 15
rect -320 -10 -252 -6
rect -245 13 -236 17
rect -212 13 -202 17
rect -245 -3 -241 13
rect -212 6 -209 13
rect -216 1 -214 5
rect -209 1 -202 5
rect -245 -7 -236 -3
rect -178 -3 -174 21
rect -297 -14 -293 -10
rect -269 -14 -265 -10
rect -464 -44 -457 -41
rect -542 -46 -511 -45
rect -461 -48 -457 -44
rect -450 -45 -437 -41
rect -429 -43 -352 -40
rect -347 -40 -309 -39
rect -347 -41 -303 -40
rect -347 -43 -296 -41
rect -564 -55 -508 -51
rect -503 -55 -498 -51
rect -652 -58 -620 -55
rect -652 -62 -649 -58
rect -671 -73 -667 -64
rect -623 -69 -620 -58
rect -550 -59 -546 -55
rect -529 -59 -525 -55
rect -508 -59 -504 -55
rect -623 -72 -577 -69
rect -749 -94 -746 -76
rect -712 -79 -583 -76
rect -696 -87 -693 -79
rect -649 -80 -583 -79
rect -635 -84 -631 -80
rect -614 -84 -610 -80
rect -593 -84 -589 -80
rect -742 -91 -655 -87
rect -756 -97 -746 -94
rect -728 -95 -724 -91
rect -707 -95 -703 -91
rect -686 -95 -682 -91
rect -665 -95 -661 -91
rect -836 -103 -813 -100
rect -817 -106 -813 -103
rect -817 -110 -809 -106
rect -782 -107 -778 -105
rect -750 -106 -746 -97
rect -817 -134 -813 -110
rect -755 -110 -746 -106
rect -750 -111 -746 -110
rect -789 -118 -779 -114
rect -755 -118 -746 -114
rect -782 -126 -779 -118
rect -789 -130 -775 -126
rect -817 -138 -809 -134
rect -750 -134 -746 -118
rect -580 -102 -577 -72
rect -574 -87 -571 -63
rect -481 -73 -477 -68
rect -483 -77 -477 -73
rect -429 -49 -426 -43
rect -473 -71 -469 -68
rect -453 -71 -449 -68
rect -473 -74 -449 -71
rect -446 -52 -426 -49
rect -446 -77 -443 -52
rect -423 -71 -420 -43
rect -306 -44 -296 -43
rect -289 -44 -285 -34
rect -277 -41 -273 -34
rect -213 -41 -209 -6
rect -182 -7 -178 -3
rect -178 -13 -174 -8
rect -280 -44 -273 -41
rect -380 -51 -325 -48
rect -277 -48 -273 -44
rect -266 -45 -262 -41
rect -169 -42 -166 146
rect -158 136 -154 166
rect -102 166 -93 170
rect -140 158 -122 162
rect -134 151 -130 158
rect -97 151 -93 166
rect -139 148 -118 151
rect -158 132 -150 136
rect -143 129 -139 146
rect -122 139 -118 148
rect -111 147 -93 151
rect -151 115 -147 119
rect -114 115 -110 119
rect -151 111 -135 115
rect -130 111 -104 115
rect -142 101 -109 105
rect -103 101 -79 105
rect -142 -3 -138 101
rect -127 97 -123 101
rect -89 97 -85 101
rect -119 70 -115 77
rect -97 70 -93 77
rect -130 66 -126 70
rect -119 66 -110 70
rect -105 66 -93 70
rect -86 66 -82 70
rect -127 40 -123 43
rect -126 35 -123 40
rect -119 37 -115 43
rect -110 45 -105 65
rect -97 63 -93 66
rect -89 37 -85 43
rect -131 20 -127 35
rect -119 34 -85 37
rect -127 15 -123 19
rect -110 18 -106 26
rect -74 19 -70 25
rect -78 15 -70 19
rect -113 7 -98 11
rect -110 2 -106 7
rect -74 -6 -70 15
rect -138 -8 -70 -6
rect -142 -10 -70 -8
rect -115 -14 -111 -10
rect -87 -14 -83 -10
rect -169 -45 -114 -42
rect -107 -44 -103 -34
rect -95 -41 -91 -34
rect -98 -44 -91 -41
rect -320 -51 -314 -48
rect -380 -52 -314 -51
rect -366 -56 -362 -52
rect -345 -56 -341 -52
rect -324 -56 -320 -52
rect -297 -73 -293 -68
rect -558 -86 -554 -79
rect -537 -86 -533 -79
rect -516 -86 -512 -79
rect -474 -80 -443 -77
rect -474 -81 -471 -80
rect -491 -84 -471 -81
rect -374 -83 -370 -76
rect -353 -83 -349 -76
rect -332 -83 -328 -76
rect -299 -77 -293 -73
rect -289 -73 -285 -68
rect -269 -73 -265 -68
rect -289 -77 -265 -73
rect -491 -86 -488 -84
rect -574 -90 -559 -87
rect -500 -90 -488 -86
rect -479 -90 -439 -87
rect -558 -94 -554 -91
rect -643 -111 -639 -104
rect -622 -111 -618 -104
rect -601 -111 -597 -104
rect -580 -105 -567 -102
rect -736 -122 -732 -115
rect -715 -122 -711 -115
rect -694 -122 -690 -115
rect -673 -122 -669 -115
rect -643 -119 -639 -116
rect -817 -144 -813 -138
rect -782 -141 -778 -137
rect -755 -138 -746 -134
rect -736 -130 -732 -127
rect -728 -171 -724 -170
rect -715 -171 -711 -170
rect -728 -174 -711 -171
rect -707 -171 -703 -170
rect -694 -171 -690 -170
rect -707 -174 -690 -171
rect -686 -171 -682 -170
rect -673 -171 -669 -170
rect -686 -174 -669 -171
rect -635 -150 -631 -149
rect -622 -150 -618 -149
rect -635 -153 -618 -150
rect -614 -150 -610 -149
rect -601 -150 -597 -149
rect -614 -153 -597 -150
rect -567 -123 -564 -105
rect -550 -125 -546 -124
rect -537 -125 -533 -124
rect -550 -128 -533 -125
rect -529 -125 -525 -124
rect -516 -125 -512 -124
rect -529 -128 -512 -125
rect -508 -125 -504 -124
rect -593 -154 -589 -149
rect -507 -154 -504 -130
rect -593 -156 -504 -154
rect -665 -171 -661 -170
rect -658 -157 -504 -156
rect -658 -159 -590 -157
rect -658 -171 -655 -159
rect -665 -174 -655 -171
rect -639 -170 -636 -159
rect -479 -160 -476 -90
rect -473 -91 -439 -90
rect -434 -91 -386 -87
rect -304 -84 -301 -78
rect -313 -87 -301 -84
rect -374 -91 -370 -88
rect -313 -91 -310 -87
rect -459 -95 -455 -91
rect -438 -95 -434 -91
rect -417 -95 -413 -91
rect -396 -95 -392 -91
rect -467 -122 -463 -115
rect -446 -122 -442 -115
rect -425 -122 -421 -115
rect -404 -122 -400 -115
rect -366 -122 -362 -121
rect -353 -122 -349 -121
rect -388 -127 -373 -124
rect -366 -125 -349 -122
rect -345 -122 -341 -121
rect -332 -122 -328 -121
rect -345 -125 -328 -122
rect -324 -122 -320 -121
rect -317 -94 -310 -91
rect -317 -122 -314 -94
rect -262 -97 -259 -46
rect -252 -105 -249 -53
rect -169 -57 -166 -45
rect -95 -48 -91 -44
rect -84 -45 -71 -41
rect -115 -73 -111 -68
rect -117 -77 -111 -73
rect -107 -73 -103 -68
rect -87 -73 -83 -68
rect -107 -77 -83 -73
rect -324 -125 -314 -122
rect -311 -108 -249 -105
rect -572 -163 -476 -160
rect -467 -130 -463 -127
rect -611 -167 -603 -164
rect -639 -174 -630 -170
rect -607 -171 -603 -167
rect -572 -170 -568 -163
rect -576 -174 -568 -170
rect -639 -182 -630 -178
rect -606 -181 -596 -178
rect -639 -200 -635 -182
rect -606 -184 -603 -181
rect -606 -192 -603 -189
rect -610 -196 -596 -192
rect -639 -204 -630 -200
rect -572 -200 -568 -174
rect -606 -213 -603 -203
rect -576 -204 -568 -200
rect -572 -210 -568 -204
rect -565 -169 -470 -166
rect -565 -213 -562 -169
rect -473 -179 -470 -169
rect -459 -171 -455 -170
rect -446 -171 -442 -170
rect -459 -174 -442 -171
rect -438 -171 -434 -170
rect -425 -171 -421 -170
rect -438 -174 -421 -171
rect -417 -171 -413 -170
rect -404 -171 -400 -170
rect -417 -174 -400 -171
rect -396 -171 -392 -170
rect -385 -179 -382 -127
rect -376 -128 -373 -127
rect -311 -128 -308 -108
rect -376 -131 -308 -128
rect -473 -182 -382 -179
rect -606 -216 -562 -213
<< metal2 >>
rect -635 202 -620 207
rect -783 185 -754 190
rect -759 163 -754 185
rect -750 127 -745 185
rect -708 158 -687 163
rect -678 127 -673 185
rect -749 117 -746 122
rect -725 119 -682 122
rect -725 117 -722 119
rect -749 114 -722 117
rect -776 92 -698 97
rect -780 77 -777 92
rect -823 74 -777 77
rect -823 -3 -820 74
rect -806 52 -803 63
rect -809 49 -803 52
rect -809 36 -806 49
rect -777 48 -704 51
rect -777 44 -774 48
rect -749 44 -746 48
rect -728 44 -725 48
rect -707 44 -704 48
rect -809 33 -803 36
rect -853 -6 -820 -3
rect -868 -72 -864 -50
rect -853 -63 -850 -6
rect -806 -7 -803 33
rect -756 5 -753 39
rect -756 2 -739 5
rect -742 -4 -739 2
rect -735 3 -732 39
rect -714 3 -711 39
rect -735 0 -718 3
rect -714 0 -689 3
rect -721 -4 -718 0
rect -742 -7 -725 -4
rect -721 -7 -696 -4
rect -815 -10 -803 -7
rect -815 -45 -812 -10
rect -728 -11 -725 -7
rect -728 -14 -703 -11
rect -706 -22 -703 -14
rect -699 -15 -696 -7
rect -692 -8 -689 0
rect -685 -1 -682 119
rect -678 82 -673 122
rect -625 82 -620 202
rect -458 190 -443 195
rect -274 190 -259 195
rect -92 190 -77 195
rect -606 173 -577 178
rect -582 151 -577 173
rect -573 115 -568 173
rect -531 146 -510 151
rect -501 115 -496 173
rect -652 68 -649 77
rect -501 70 -496 110
rect -448 70 -443 190
rect -422 173 -393 178
rect -398 151 -393 173
rect -389 115 -384 173
rect -347 146 -326 151
rect -317 115 -312 173
rect -317 70 -312 110
rect -264 70 -259 190
rect -240 173 -211 178
rect -216 151 -211 173
rect -207 115 -202 173
rect -165 146 -144 151
rect -135 115 -130 173
rect -135 70 -130 110
rect -82 70 -77 190
rect -568 56 -427 61
rect -384 56 -245 61
rect -202 56 -61 61
rect -476 31 -471 40
rect -523 26 -476 29
rect -647 4 -579 7
rect -647 0 -644 4
rect -624 0 -621 4
rect -603 0 -600 4
rect -582 0 -579 4
rect -523 0 -520 26
rect -430 8 -427 56
rect -412 31 -332 34
rect -292 31 -287 40
rect -412 8 -409 31
rect -295 27 -292 29
rect -370 24 -292 27
rect -402 12 -379 15
rect -402 8 -399 12
rect -382 8 -379 12
rect -370 8 -367 24
rect -342 8 -293 11
rect -430 5 -425 8
rect -685 -4 -647 -1
rect -557 -4 -520 0
rect -481 -3 -477 2
rect -424 -1 -420 3
rect -403 -1 -399 3
rect -424 -4 -399 -1
rect -692 -9 -652 -8
rect -692 -11 -655 -9
rect -634 -11 -631 -5
rect -634 -14 -627 -11
rect -699 -18 -660 -15
rect -706 -25 -667 -22
rect -663 -23 -660 -18
rect -670 -29 -667 -25
rect -794 -34 -717 -31
rect -670 -32 -647 -29
rect -794 -45 -791 -34
rect -785 -41 -761 -38
rect -785 -45 -782 -41
rect -764 -45 -761 -41
rect -720 -43 -717 -34
rect -663 -41 -659 -36
rect -841 -49 -828 -46
rect -827 -54 -824 -50
rect -806 -54 -803 -50
rect -785 -54 -782 -50
rect -827 -57 -782 -54
rect -868 -75 -811 -72
rect -814 -97 -811 -75
rect -814 -100 -780 -97
rect -773 -98 -770 -50
rect -705 -81 -702 -41
rect -650 -46 -647 -32
rect -652 -49 -647 -46
rect -652 -59 -649 -49
rect -630 -51 -627 -14
rect -630 -54 -618 -51
rect -652 -62 -625 -59
rect -628 -74 -625 -62
rect -621 -67 -618 -54
rect -613 -59 -610 -5
rect -592 -9 -589 -5
rect -592 -12 -521 -9
rect -524 -14 -521 -12
rect -524 -17 -465 -14
rect -519 -41 -512 -38
rect -468 -40 -465 -17
rect -613 -62 -575 -59
rect -621 -70 -571 -67
rect -628 -77 -578 -74
rect -773 -101 -742 -98
rect -745 -123 -742 -101
rect -720 -99 -717 -81
rect -705 -84 -585 -81
rect -720 -102 -700 -99
rect -736 -118 -712 -115
rect -736 -122 -733 -118
rect -715 -122 -712 -118
rect -703 -122 -700 -102
rect -694 -118 -670 -115
rect -694 -122 -691 -118
rect -673 -122 -670 -118
rect -660 -122 -657 -84
rect -643 -107 -598 -104
rect -643 -111 -640 -107
rect -622 -111 -619 -107
rect -601 -111 -598 -107
rect -588 -111 -585 -84
rect -581 -116 -578 -77
rect -574 -109 -571 -70
rect -547 -79 -544 -48
rect -515 -66 -512 -41
rect -427 -45 -394 -42
rect -427 -51 -424 -45
rect -445 -54 -424 -51
rect -515 -69 -502 -66
rect -566 -82 -544 -79
rect -566 -100 -563 -82
rect -547 -86 -544 -82
rect -536 -82 -514 -79
rect -536 -86 -533 -82
rect -517 -86 -514 -82
rect -505 -86 -502 -69
rect -445 -79 -442 -54
rect -397 -56 -394 -45
rect -404 -59 -394 -56
rect -473 -82 -442 -79
rect -493 -85 -470 -82
rect -557 -95 -554 -91
rect -538 -95 -535 -91
rect -557 -98 -535 -95
rect -524 -95 -521 -91
rect -493 -95 -490 -85
rect -524 -98 -490 -95
rect -423 -100 -420 -76
rect -397 -90 -394 -59
rect -390 -83 -387 3
rect -342 -6 -337 8
rect -248 9 -245 56
rect -110 31 -105 40
rect -208 26 -110 31
rect -248 6 -209 9
rect -327 -2 -280 1
rect -363 -43 -352 -40
rect -363 -83 -360 -43
rect -325 -46 -322 -11
rect -283 -40 -280 -2
rect -110 -27 -107 -3
rect -253 -30 -107 -27
rect -253 -41 -250 -30
rect -257 -44 -250 -41
rect -208 -44 -103 -41
rect -66 -45 -61 56
rect -314 -53 -253 -50
rect -71 -50 -66 -46
rect -248 -53 -66 -50
rect -353 -79 -328 -76
rect -353 -83 -349 -79
rect -332 -83 -328 -79
rect -314 -83 -311 -53
rect -264 -60 -170 -57
rect -264 -82 -261 -60
rect -390 -86 -375 -83
rect -397 -93 -379 -90
rect -562 -105 -452 -102
rect -574 -112 -486 -109
rect -745 -126 -737 -123
rect -777 -145 -743 -142
rect -746 -176 -743 -145
rect -723 -148 -720 -127
rect -715 -131 -712 -127
rect -694 -131 -691 -127
rect -715 -134 -691 -131
rect -681 -139 -678 -127
rect -630 -132 -627 -116
rect -611 -125 -608 -116
rect -581 -119 -550 -116
rect -611 -128 -569 -125
rect -630 -135 -579 -132
rect -681 -141 -583 -139
rect -567 -141 -564 -128
rect -553 -130 -550 -119
rect -489 -123 -486 -112
rect -455 -122 -452 -105
rect -434 -103 -420 -100
rect -382 -99 -379 -93
rect -374 -92 -370 -88
rect -354 -92 -349 -88
rect -374 -95 -349 -92
rect -316 -87 -311 -83
rect -307 -85 -261 -82
rect -342 -92 -337 -88
rect -307 -92 -304 -85
rect -342 -95 -304 -92
rect -382 -102 -264 -99
rect -434 -122 -431 -103
rect -255 -106 -252 -60
rect -310 -109 -252 -106
rect -426 -118 -400 -115
rect -426 -122 -423 -118
rect -403 -122 -400 -118
rect -489 -126 -468 -123
rect -553 -133 -514 -130
rect -517 -134 -514 -133
rect -467 -131 -464 -127
rect -446 -131 -443 -127
rect -425 -131 -422 -127
rect -467 -134 -422 -131
rect -413 -131 -410 -127
rect -310 -131 -307 -109
rect -413 -134 -307 -131
rect -517 -135 -500 -134
rect -517 -137 -472 -135
rect -503 -138 -472 -137
rect -413 -138 -410 -134
rect -475 -141 -410 -138
rect -681 -142 -564 -141
rect -586 -144 -564 -142
rect -723 -151 -540 -148
rect -746 -179 -640 -176
rect -643 -185 -640 -179
rect -643 -188 -607 -185
<< m123contact >>
rect -778 208 -773 213
rect -705 208 -700 213
rect -640 202 -635 207
rect -720 193 -715 198
rect -648 193 -643 198
rect -788 185 -783 190
rect -759 158 -754 163
rect -750 185 -745 190
rect -678 185 -673 190
rect -713 158 -708 163
rect -687 158 -682 163
rect -750 122 -745 127
rect -678 122 -673 127
rect -781 92 -776 97
rect -698 92 -693 97
rect -802 40 -797 45
rect -779 39 -774 44
rect -758 39 -753 44
rect -749 39 -744 44
rect -737 39 -732 44
rect -728 39 -723 44
rect -716 39 -711 44
rect -707 39 -702 44
rect -695 39 -690 44
rect -869 -50 -864 -45
rect -652 113 -646 118
rect -601 196 -596 201
rect -528 196 -523 201
rect -417 196 -412 201
rect -344 196 -339 201
rect -235 196 -230 201
rect -162 196 -157 201
rect -463 190 -458 195
rect -279 190 -274 195
rect -97 190 -92 195
rect -543 181 -538 186
rect -471 181 -466 186
rect -611 173 -606 178
rect -582 146 -577 151
rect -573 173 -568 178
rect -501 173 -496 178
rect -536 146 -531 151
rect -510 146 -505 151
rect -573 110 -568 115
rect -501 110 -496 115
rect -678 77 -673 82
rect -653 77 -648 82
rect -625 77 -620 82
rect -475 101 -469 106
rect -359 181 -354 186
rect -287 181 -282 186
rect -427 173 -422 178
rect -398 146 -393 151
rect -389 173 -384 178
rect -317 173 -312 178
rect -352 146 -347 151
rect -326 146 -321 151
rect -389 110 -384 115
rect -317 110 -312 115
rect -501 65 -496 70
rect -476 65 -471 70
rect -448 65 -443 70
rect -291 101 -285 106
rect -177 181 -172 186
rect -105 181 -100 186
rect -245 173 -240 178
rect -216 146 -211 151
rect -207 173 -202 178
rect -135 173 -130 178
rect -170 146 -165 151
rect -144 146 -139 151
rect -207 110 -202 115
rect -135 110 -130 115
rect -317 65 -312 70
rect -292 65 -287 70
rect -264 65 -259 70
rect -109 101 -103 106
rect -135 65 -130 70
rect -110 65 -105 70
rect -82 65 -77 70
rect -573 56 -568 61
rect -389 56 -384 61
rect -207 56 -202 61
rect -674 45 -669 50
rect -476 40 -471 45
rect -497 35 -492 40
rect -476 26 -471 31
rect -498 15 -493 20
rect -368 39 -363 44
rect -325 40 -320 45
rect -292 40 -287 45
rect -332 31 -327 36
rect -313 33 -308 38
rect -292 26 -287 31
rect -314 15 -309 20
rect -425 3 -420 8
rect -413 3 -408 8
rect -404 3 -399 8
rect -392 3 -387 8
rect -383 3 -378 8
rect -371 3 -366 8
rect -647 -5 -642 0
rect -635 -5 -630 0
rect -626 -5 -621 0
rect -614 -5 -609 0
rect -605 -5 -600 0
rect -593 -5 -588 0
rect -584 -5 -579 0
rect -562 -5 -557 0
rect -477 -3 -472 2
rect -655 -14 -650 -9
rect -705 -41 -700 -36
rect -684 -41 -679 -36
rect -668 -41 -663 -36
rect -846 -50 -841 -45
rect -828 -50 -823 -45
rect -816 -50 -811 -45
rect -807 -50 -802 -45
rect -795 -50 -790 -45
rect -786 -50 -781 -45
rect -774 -50 -769 -45
rect -765 -50 -760 -45
rect -721 -48 -716 -43
rect -853 -68 -848 -63
rect -748 -58 -743 -53
rect -749 -76 -744 -71
rect -667 -73 -662 -68
rect -508 -10 -503 -5
rect -448 -10 -443 -5
rect -547 -48 -542 -43
rect -575 -54 -570 -49
rect -575 -63 -570 -58
rect -783 -105 -778 -100
rect -644 -116 -639 -111
rect -632 -116 -627 -111
rect -623 -116 -618 -111
rect -611 -116 -606 -111
rect -602 -116 -597 -111
rect -590 -116 -585 -111
rect -469 -45 -464 -40
rect -437 -46 -432 -41
rect -508 -55 -503 -50
rect -488 -78 -483 -73
rect -424 -76 -419 -71
rect -559 -91 -554 -86
rect -547 -91 -542 -86
rect -538 -91 -533 -86
rect -526 -91 -521 -86
rect -517 -91 -512 -86
rect -505 -91 -500 -86
rect -439 -91 -434 -86
rect -293 6 -288 11
rect -110 40 -105 45
rect -131 35 -126 40
rect -213 26 -208 31
rect -110 26 -105 31
rect -241 21 -236 26
rect -132 15 -127 20
rect -332 -2 -327 3
rect -214 1 -209 6
rect -342 -11 -337 -6
rect -325 -11 -320 -6
rect -374 -36 -369 -31
rect -352 -43 -347 -38
rect -111 -3 -106 2
rect -178 -8 -173 -3
rect -143 -8 -138 -3
rect -285 -45 -280 -40
rect -262 -46 -257 -41
rect -213 -46 -208 -41
rect -103 -45 -98 -40
rect -71 -46 -66 -41
rect -325 -51 -320 -46
rect -253 -53 -248 -48
rect -304 -78 -299 -73
rect -375 -88 -370 -83
rect -363 -88 -358 -83
rect -354 -88 -349 -83
rect -567 -105 -562 -100
rect -737 -127 -732 -122
rect -725 -127 -720 -122
rect -716 -127 -711 -122
rect -704 -127 -699 -122
rect -695 -127 -690 -122
rect -683 -127 -678 -122
rect -674 -127 -669 -122
rect -662 -127 -657 -122
rect -782 -146 -777 -141
rect -569 -128 -564 -123
rect -342 -88 -337 -83
rect -333 -88 -328 -83
rect -321 -88 -316 -83
rect -264 -102 -259 -97
rect -170 -62 -165 -57
rect -122 -78 -117 -73
rect -508 -130 -503 -125
rect -468 -127 -463 -122
rect -456 -127 -451 -122
rect -447 -127 -442 -122
rect -435 -127 -430 -122
rect -426 -127 -421 -122
rect -414 -127 -409 -122
rect -405 -127 -400 -122
rect -393 -127 -388 -122
rect -616 -167 -611 -162
rect -396 -176 -391 -171
rect -607 -189 -602 -184
<< metal3 >>
rect -681 226 -595 230
rect -773 208 -705 213
rect -778 114 -773 208
rect -681 198 -676 226
rect -598 218 -595 226
rect -598 215 -133 218
rect -598 214 -315 215
rect -715 194 -648 198
rect -652 193 -648 194
rect -596 196 -528 201
rect -652 118 -646 193
rect -778 111 -682 114
rect -698 97 -695 111
rect -685 92 -682 111
rect -601 92 -596 196
rect -504 186 -499 214
rect -412 196 -344 201
rect -538 182 -471 186
rect -475 181 -471 182
rect -475 106 -469 181
rect -417 92 -412 196
rect -320 186 -315 214
rect -230 196 -162 201
rect -354 182 -287 186
rect -291 181 -287 182
rect -291 106 -285 181
rect -235 92 -230 196
rect -138 186 -133 215
rect -172 182 -105 186
rect -109 181 -105 182
rect -109 106 -103 181
rect -685 89 -230 92
rect -685 50 -682 89
rect -685 46 -674 50
rect -811 41 -802 44
rect -811 -6 -808 41
rect -693 5 -690 39
rect -601 40 -596 89
rect -417 52 -412 89
rect -417 49 -310 52
rect -601 36 -497 40
rect -836 -9 -808 -6
rect -705 2 -690 5
rect -836 -56 -833 -9
rect -705 -36 -702 2
rect -683 -45 -680 -41
rect -716 -48 -680 -45
rect -756 -56 -748 -53
rect -836 -59 -766 -56
rect -769 -99 -766 -59
rect -769 -102 -760 -99
rect -763 -119 -760 -102
rect -756 -112 -753 -56
rect -665 -54 -575 -51
rect -570 -54 -567 36
rect -363 40 -325 44
rect -363 39 -347 40
rect -313 38 -310 49
rect -235 40 -230 89
rect -235 36 -131 40
rect -235 26 -230 36
rect -236 21 -230 26
rect -508 -50 -505 -10
rect -665 -68 -662 -54
rect -736 -71 -667 -68
rect -736 -72 -733 -71
rect -744 -75 -733 -72
rect -496 -73 -493 15
rect -496 -77 -488 -73
rect -756 -115 -644 -112
rect -763 -122 -741 -119
rect -744 -152 -741 -122
rect -496 -125 -493 -77
rect -446 -83 -443 -10
rect -435 -11 -342 -8
rect -435 -41 -432 -11
rect -313 -31 -309 15
rect -173 -7 -143 -3
rect -369 -34 -309 -31
rect -437 -58 -434 -46
rect -313 -73 -309 -34
rect -131 -73 -127 15
rect -313 -77 -304 -73
rect -131 -77 -122 -73
rect -446 -86 -434 -83
rect -503 -128 -493 -125
rect -497 -132 -493 -128
rect -497 -135 -393 -132
rect -744 -155 -611 -152
rect -614 -162 -611 -155
rect -396 -171 -393 -135
<< m234contact >>
rect -806 63 -801 68
rect -653 63 -648 68
rect -660 -25 -655 -20
rect -659 -41 -654 -36
rect -524 -41 -519 -36
rect -486 -3 -481 2
rect -721 -81 -716 -76
rect -438 -63 -433 -58
rect -409 -60 -404 -55
rect -579 -137 -574 -132
rect -540 -152 -535 -147
<< metal4 >>
rect -801 64 -653 67
rect -667 12 -502 15
rect -667 -29 -664 12
rect -505 2 -502 12
rect -505 -1 -486 2
rect -655 -23 -531 -20
rect -667 -32 -656 -29
rect -659 -36 -656 -32
rect -650 -77 -647 -23
rect -534 -26 -531 -23
rect -534 -29 -521 -26
rect -524 -36 -521 -29
rect -408 -55 -405 -51
rect -437 -67 -434 -63
rect -716 -80 -647 -77
rect -578 -70 -434 -67
rect -578 -132 -575 -70
rect -408 -96 -405 -60
rect -539 -99 -405 -96
rect -539 -147 -536 -99
<< labels >>
rlabel metal3 -138 214 -133 218 1 vdd
rlabel m123contact -170 146 -165 151 1 p_0
rlabel metal1 -110 1 -106 5 1 g_0
rlabel m123contact -135 110 -130 115 1 b_0
rlabel metal2 -82 143 -77 148 1 a_0
rlabel m123contact -207 110 -202 115 1 c0
rlabel m123contact -245 173 -240 178 1 s0
rlabel metal3 -235 36 -230 40 1 gnd
rlabel m123contact -427 173 -422 178 3 s1
rlabel m123contact -352 146 -347 151 1 p_1
rlabel m123contact -389 110 -384 115 1 c1
rlabel m123contact -317 110 -312 115 1 b_1
rlabel metal2 -264 143 -259 148 1 a_1
rlabel metal1 -102 -44 -97 -41 1 p0c0
rlabel m123contact -292 26 -287 31 1 gb_1
rlabel m123contact -110 26 -105 31 1 gb_0
rlabel metal1 -284 -44 -279 -41 1 p1g0
rlabel m123contact -375 -88 -370 -83 1 p1p0c0
rlabel m123contact -573 110 -568 115 1 c2
rlabel metal2 -448 143 -443 148 1 a_2
rlabel m123contact -501 110 -496 115 1 b_2
rlabel m123contact -536 146 -531 151 1 p_2
rlabel metal1 -476 1 -472 5 1 g_2
rlabel m123contact -476 26 -471 31 1 gb_2
rlabel metal1 -468 -44 -463 -41 1 p2g1
rlabel m123contact -611 173 -606 178 3 s2
rlabel m123contact -559 -91 -554 -86 1 p2p1g0
rlabel metal3 -468 -127 -463 -122 1 p2p1p0c0
rlabel metal2 -625 145 -620 150 1 a_3
rlabel m123contact -678 122 -673 127 1 b_3
rlabel m123contact -788 185 -783 190 3 s3
rlabel m123contact -293 6 -288 11 1 g_1
rlabel m123contact -697 94 -695 95 1 gnd
rlabel metal1 -668 -72 -664 -70 8 gnd
rlabel m123contact -704 -40 -701 -37 1 p_3
rlabel metal1 -688 -40 -684 -38 1 p3g2
rlabel metal1 -555 -53 -552 -52 1 vdd
rlabel metal1 -686 -5 -686 -5 1 vdd
rlabel metal1 -590 -157 -586 -156 8 gnd
rlabel m123contact -567 -105 -562 -100 1 p_2
rlabel metal1 -620 -79 -619 -78 1 vdd
rlabel polycontact -594 -115 -590 -111 1 p_3
rlabel m123contact -644 -116 -639 -111 1 p3p2g1
rlabel metal1 -689 -89 -685 -88 5 vdd
rlabel polycontact -687 -126 -683 -122 1 p_2
rlabel polycontact -708 -126 -704 -122 1 p_1
rlabel polycontact -530 -90 -526 -86 1 g_0
rlabel m123contact -737 -127 -732 -122 1 p3p2p1g0
rlabel metal1 -783 6 -783 6 1 vdd
rlabel metal1 -787 -12 -787 -12 1 vdd
rlabel metal1 -753 -96 -753 -96 1 gnd
rlabel metal1 -796 41 -796 41 1 p
rlabel metal1 -638 -171 -636 -167 4 gnd
rlabel metal1 -606 -191 -604 -187 3 out
rlabel metal1 -570 -180 -570 -180 1 vdd
rlabel metal1 -607 -170 -603 -165 1 p
rlabel metal1 -749 -107 -747 -103 6 gnd
rlabel metal1 -815 -131 -813 -118 3 vdd
rlabel metal1 -606 -210 -603 -204 1 c0
rlabel metal1 -781 -129 -779 -127 1 c4
rlabel m123contact -647 -5 -642 0 1 c3
rlabel m123contact -562 -5 -557 0 1 gb_2
rlabel m123contact -713 158 -708 163 1 p_3
rlabel m123contact -652 79 -652 79 1 gb_3
rlabel metal1 -866 -10 -866 -10 4 vdd
rlabel m123contact -781 -103 -781 -103 1 gb
rlabel m123contact -828 -50 -823 -45 1 g
<< end >>
