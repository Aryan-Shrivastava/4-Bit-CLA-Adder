.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={10*LAMBDA}
.param width_P={20*LAMBDA}
.global gnd vdd

Vdd	vdd	gnd	'SUPPLY'
va x gnd pulse (0 1.8 0 0.1n 0.1n 1n 2n)
*******************************************************************************************************************************************************
* Inverter Circuit
.subckt inv y x vdd gnd 
    M1 y x gnd gnd  CMOSN W={width_N} L={2*LAMBDA} AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    M2 y x vdd vdd  CMOSP W={width_P} L={2*LAMBDA} AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv
xinv y x vdd gnd inv
.tran 0.1n 20n

.control
set color0=white
run 
plot v(x) v(y)+2
.endc