magic
tech scmos
timestamp 1731333581
<< nwell >>
rect -84 47 -22 81
<< ntransistor >>
rect -73 8 -71 38
rect -54 8 -52 38
rect -35 8 -33 38
<< ptransistor >>
rect -73 53 -71 73
rect -54 53 -52 73
rect -35 53 -33 73
<< ndiffusion >>
rect -74 8 -73 38
rect -71 8 -70 38
rect -55 8 -54 38
rect -52 8 -51 38
rect -36 8 -35 38
rect -33 8 -32 38
<< pdiffusion >>
rect -74 53 -73 73
rect -71 53 -70 73
rect -55 53 -54 73
rect -52 53 -51 73
rect -36 53 -35 73
rect -33 53 -32 73
<< ndcontact >>
rect -78 8 -74 38
rect -70 8 -66 38
rect -59 8 -55 38
rect -51 8 -47 38
rect -40 8 -36 38
rect -32 8 -28 38
<< pdcontact >>
rect -78 53 -74 73
rect -70 53 -66 73
rect -59 53 -55 73
rect -51 53 -47 73
rect -40 53 -36 73
rect -32 53 -28 73
<< polysilicon >>
rect -73 73 -71 76
rect -54 73 -52 76
rect -35 73 -33 76
rect -73 38 -71 53
rect -54 38 -52 53
rect -35 38 -33 53
rect -73 4 -71 8
rect -54 4 -52 8
rect -35 4 -33 8
<< polycontact >>
rect -77 42 -73 46
rect -58 42 -54 46
rect -39 42 -35 46
<< metal1 >>
rect -84 77 -22 81
rect -78 73 -74 77
rect -59 73 -55 77
rect -40 73 -36 77
rect -70 46 -66 53
rect -51 46 -47 53
rect -32 46 -28 53
rect -32 38 -28 41
rect -78 3 -74 8
rect -82 -1 -74 3
rect -70 3 -66 8
rect -59 3 -55 8
rect -70 -1 -55 3
rect -51 3 -47 8
rect -40 3 -36 8
rect -51 -1 -36 3
<< metal2 >>
rect -65 41 -51 46
rect -46 41 -32 46
<< m123contact >>
rect -70 41 -65 46
rect -51 41 -46 46
rect -32 41 -27 46
<< labels >>
rlabel metal1 -81 0 -77 1 2 gnd
rlabel metal1 -56 79 -52 80 5 vdd
rlabel polycontact -77 42 -73 46 1 a
rlabel polycontact -58 42 -54 46 1 b
rlabel polycontact -39 42 -35 46 1 c
rlabel m123contact -32 41 -27 46 1 out
<< end >>
